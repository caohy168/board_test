`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
jXsoZcqMe6B1UnGf9hyp9ifP9jk4P+1XJJAI0ZVRLEzDYWGbO1NPI0RDqIVdaf9s7Vr5j9uazwKz
Ns/gABC7FA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
if7S2GOcV3J9rYyUQpwBUXgCuzD4IEfYkh9IFRilZAgECja0nXBOBfZZG6c4L6vtGmj9Yzq71wZd
Xlk2LkjFCvg7RkmgORflZy2j/Sz7D5ft8xyiRpirF87XLe87AdPJVNS4hLsnkffkAxfZo4yyF0Fj
yGP4cfAaVIUtXGb61hg=

`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
C4JYOuQq5u95wgv01rUHguZ95v+CjaL+kVpziQFbJ4BXjYg6pORftttbleiVh7aJ+3Ct8xOWcHnB
vIdiwDM3LZigPzxYXFAXpnV3wxg0k+q6OWfmi1a9lnEDB1eIqxTWvy+0z3TbQhhWbuE4/A5KapYD
0TZHB0Hyi/x+1faZd88=

`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
xhKhbS2zpuVWlO6/Qj5Lj7VDSzriDCw//I3BIyThxOPBYxOwYenXNCb18Slf5Eq7Ca4ooPTljSWz
rkstZtGXwjjGrnfK08ibqtJ+epHFsv2HrCa9EejWWeytlnyMD4LTfSKLfUe43c83iQ14e3p+2LyL
FGod2Lq6Qpw6J8Sz+BbyRsA850Z8jvVtSsSApvGv3aPIzKZkU52aMTPwjsmGj82XOMpNjbMAft7n
LSASdR1aSzWh14gLc1mrCjzJMQo6PNsejUkv5dsPeLgWqUtVjAnGlbDhml8kRPHza99S8ZUL+WuM
25Kd4o6yKILqaEZ3XTEmNh4aw+GbR9JGzDd+Dg==

`pragma protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
IV3N1NDZDtplL6tSmUZLRIqyEFSv3B+hsLg6K1ngz6C2q6IDEx9mrrsfad1gbSxx+DSxVQIWrRGw
tK8ADcuK4oYCPF5BLDhAriZbOja4zvyaufPcfwub60hOlMTzu2ZBJ0Gcj36WazzpMEwwahIuTER3
oFD02d1tCg2QP61RQssnC2Rq/U4vvpim4KMuqPVnS8V6YdLZqYAo/za/1H4vm4XhrAWtd/XrmXD3
yHI13YSuJBbyNvGodALO/LLQNEzsCqaxZxh6MvPWDi34NckHU17XutUcIBxgbie3B1kejcs8f6t+
CcjwtDOZnjxYfLAAgs4gDbfx1g2tYBCSlagJCQ==

`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
DEfZcZQ3VHU29kiHHkCcusZNaoJ1kx6jQnIMklaa+bRtmwTH9LQTiki+e3u9c5SHYMd769t2xCWp
LMLv8nNuAIgzaQLSx+JRNzhPpynFsA6EKsJLX3j/3ilurljgloAOIb5+LvX9jWtYSrq3RxZrHFkZ
cRSOcA8XeNVWIRoJcHDDsvRwFdTuxSXCN4ikJ0FMvQ7kS912pDYaG1HSZgiVgbQwJLhF/+X/axl7
nAwsknFCkOmWSJyAQE85vLAlKegt58FtS4zdtplpOOl4QXpBEUBxWyztHxDLz5C2U/KPeudxasq+
EPg7zp5LpKU/M9m/UE5ETCrTnC7NxkfwVjeOiQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 827600)
`pragma protect data_block
4bLjqS4aA4KqhBmAjPx/dTxidPbtPaUeBP8+jxvxQU12iK0YVXpnRAZ7kF5W26vPIV06u7FzInpA
li9JUFnxhAl7O9LAktlfIWQjDjnKenvCDi9vVXsnXA6QYLxBu0mDxu1Fnu+jUup3hEpKuhkPy+bH
3qzR89NX5wXLfCVAfycBV7sX5kO7Fe3ecrnlBOOs2kYZtWM0cPSJzFP1VF9Az9sUYDNwGy2D+0Or
b9+q3xoSuIRfQzQiOAdUI9BZxExxcpDiMiX0ZGwT8HhoV+n+JDaCOUZO6r/MB3FYFrB8Y+JaW3FO
xgVenFkrYkjSyv7JN2D86wDxdK3wC+tXd8H5MngXzM2+X4H+8cbCHi3S0GgwLB/yR1aGs8/rtjQ6
e82N6Aotwfka64ucBywgrCLFloz8xr8HvLI6PCpsLrCFcG5RA3BJEODB79CO+0TU/J5vec0Y5nQ9
EDhqiPSopQGzv3RTCNuduKj5Mi1BhGhREigJrxjQzmG+no9YBOyMKb+T0DA8TFB8Ht2CiqfqsYWG
k2f2MjaR7bBKtxT4CwmbesUo99qU75QimMQBOKW+rY3omze1veJ42P2egFV71J+UveXvez5W+ag7
rKAsZNLgRITMRgH4HVgw94RK0lNB8mqKfgwCfxk5MW9vqC3vxe7WL7FHO52owmmXEjnxWGaI6bQW
skyXvPfQZ8Su9uvVo0rReI7V+WSbZvzrTG2Gu2nXCIYaf1RfJFDZSit49SdCCXG37b4oOxQmv8zW
CB1t8zxTmePj9DM3GSFLZs/DP+jfG8kCCCe/D8Dzvh2x9Rxr9/HbG/yMDlBI7+S/7qbB6NYe1rVh
dWgn2+HDN41JcsJgn2hG0lbc6B4rGDUvURaUExKO2nHZM7Q20OUeZRst9nW6cVEl6bQDetv6TvVH
IQeWDWjFM6bHKkPH5mvqG1gtLsOah6rLiJk9Dn5dAcur4ZyfE5JCkZRdjlQc0Kwclmfx59vTTITN
32DJeNPoVU18376AB3QeNC8Yu6Jv6ZWMGxL0sRPrD1B1c89vZolMNIgBlCrSynbAXysc7J7eN6EF
94rGzGp0eRpdz6mS8LW26SY+Jc+/AwO11GEEkBaWAlgec6JsIhyJn+QjlG3FoQhmIWCKwRqZd24P
z2ktq7Ds9NT2Sr2OdpPzvxyhVnb5P0CcYAEqvm76dx8GFlWpJTbt4Vp0msHP8UrJRFkkzEXiUs8X
xqD5FWaSzQOI0g0b1jjxqmmTi5H2FzBDWWckYQBwUV5EfD/rTMiFjy4GuTOIBoJxQZW0v9NWgoxC
AnjOXOqP0K4wvddPx5kxv8wRWSmCZZtO1Lsu9OZc6zDPH0FsJHuNUwNrO/zx3komKbeZTjkKAx+q
3cDgujXJdU1eP6SsSlq23CeP9GxeXaxode4uh8oqOCZ050W1ItZf0FLdiXwCz9pTBICqwXUQsJ8+
6QlHlz+xPbWOG4BkmHafDi6YLSuNjKohLBxD2AuFAVQzKJLXlXEbq3Cmgx5UzfZR4tMVo3dJHbtV
4cbDHpKfEgz8ghw5JlpOw122Fa8zomDZCnwt79lVTaw6zJHiNduM4KEma0fnh2Ea2R5DzfjlS67l
SwFcMl8awI7ka1Bu3pBJF5r8cdMfvj+GxPBgPCGDfP/vIoxa44xAoPE0S9ozl1dWGyT3zZbzOtge
hkP+4Af6rqzPULyVumHl46ZqFCVdASz0JtvFYd934aPWSeXbXOAu2QEsnqHKa1ly5ZwHgk3q/riM
viYg6V0Tjukf8npDzDXneamSgZ8ADT7wPgNk+3t28gKIcNFcFN9oYeBMQ8etjTAiQpGBK/F7m0mD
5bf2Cl7ytNyce/ObvlWv0pGakFIP8B1euduLy4igZ+9ny+BHtwElOKzfQL4Zta1I6Cr4dsKa4OVJ
nK0P/OphtPz1C5In5++3NrVpyhw3amaBoVvCESaElBjF8YOj3kGU2ysDj0fFDfUWJOVDlvSSMzIc
N8X56DiUpnJb5LxuVYAbyyX7Po815nM4ylSAd7I+uWp/xUbjgGhE8hnh/lCpjZhzUzJTopt0UuzK
0aq6V5f2U5J4i53bo83qpCt7Tvqt0n/Tb/IgCJ7ciK9acgknkxbwWHHGphw4rp8Kyk6r3rId259Z
u+DMWhUeiNpoK0qBiYZ/NQHh/ZJADHCD3WuguEDkEcYRuyYIhJ4KzKzT4Cl2bpHl/Nd/rF2a/avN
l6JE56SmJW73qrHEsOJqurtcu4f7DoUsdGNgaMkdkjMA8GXC03cQYmLTZqYu+JAqpgui6qV5ntNu
tCsJWXNLHQFvCMvn8/2pvtHeL8kFtLA/YK64Nyp23NgF9bu8oeA6VQsNNuoQbVJygHNe2Wo1JejR
YmyIIWxCH+GTv98+w3eSHCn9u/oduzXRAInpwg6813o9cX+/g/tvh6H2X1EWLh1v5IQk0y2Ky07R
hLoI2MSmt1WrMGWvipcDjAscMDzumzGz6P4O2Ls5ZzMDGHpZHZTxz3R7wJBnXloLNDDoedEysc1P
fAGZkvKSeFlegyj8ignDwlii3RDLiJ2yEP9TERUZQds36lkEwJmP/hW/JUqHcs2WfVZEnub+Ubs7
gK5F9DPPpzYerXnI0HzL1PV7jCp9flPDZuw97KxqkzwVZ/PeHhKWJo6F+Q8A3LWQZSw3LKHOSPWj
qoVSMoaSgpyXPM5RmFm+CENWHuDLPBe/MDVfA3NIpDyQhEsJIo8elaL/1c26okBhKfaTDHJ8wzig
miwFdGWTQJg4Ez/pGc7f5S/99l1UihvB+5A6pnN2YOvw8WwSdmv827tu8dy8YCU3xRkK9SPIh6Hc
JZqn2OOguCGtIhJibvEBFNwMOX99QMlKDeNWoydg/UqE6+1i6aNm9UJ2naYZiDgTKCkl/Tc9NEM4
JRkQD5tL/sgsfdR3kbCmwFQ4lVKZZN8CISUu7VWM4u3qPqpqZ6zKTaDx/66jx4u/zEBgOqJ3W8fM
8Rsw+Sc0NocwBLhjibcmdcBYb9TrjEFzKjNhWL77AvI+Us3iMyVdSmQ93WSa4OAzD0fOg9nn5hKV
2Yhb4CvKDj2gTbCw4bK8fDQYl8n34VuUa81D73OJr5ifRzmZIOXsO1vGP5KWb/zkslHf51rDK31V
vw846gd5G1dpNFpg744OM8WSSXMfVRtD9xVuts27+o5e9nUEiFzIQgZODC+5BxONb27g8L513um4
M+pGFgPtw/UTWArSrP1dkTXVG3lUYkuGyC42kG+2aGigkO1M+l2vGLhcmtpBOxPcluZ7Lp5APr13
Ru9LP3fPiUT9YiLr/35k60Pe5BIwP9Pxz0BmH7AP2J6Ogeur9uu8kL6AzFtKxSi7X8Xj/RP288gQ
1jA/EV5DBgiHRHhe2FQnVzlH20gDp9H397dYHWEMW6PH+DMZmTlQPhwGpMwZ8P4fA/dB6rv957eV
JI5pO1/0yw0wSxK2pj5mPxhrGeC1iLajOw9z5loZyp85kjvHYaW3b6VMfAgoH5crGYu0wNwwnxXJ
XJhpanpmnhxe8DSKkAyE7Vc6kQzQcNCVbB7evpFhRdHYxfp3VAMFp2zAoMaCcdE47EUbwioyg1Mk
6vDk7BTRxS9P6WVtVRKFuc+bzHppOcujioMWTMcFBXklWBwqi1p8JG5OARj5KmIpRcTjuQTRT3wl
ADNq8xobQ652KyVp2pxTFtD4smbKi6Iy86ALfYptwUxTDXxNX8rN71KJknJy49BkRDoBdJWE3lgF
hqN23CaB5VUzjSyPimZiyhuRBBCncQHZPQzEl9mj6o5a/dP2g5UGPIqYGg7CpJaGWNyrLY05Dioh
5zLSsIwhQ9T5VIsbmQcqRX71bAPC7Hjdl2XY6g9sNiXKqnHo9yZDnXE3PFmCLQ17CKAP0t/E2EOF
29M5AE5sPfJY6Msywt1CY/oX0YkXfr4P2ICpuDhzfWHRM/ktgvp5sY4Ya6UPQfr0VV1VzmthOySK
hAm0yexU7D82ikmIjacobJ8GTwEpXdlNWcxV8eAJO96rJZTRcR6HdqxILNqkQzxVXzzEg8Gvd24C
EO3kN8ZmM9JA2p9ueDddt2Ud5k736VvJXqWAVtmWe2fh4Y/l02Glhn3DBb6govLP+ku13HhWmXvp
maoqppKSN/hMPW0Qbj+hmXo4ompHInO2oNeOxtPmrA16/gfx6OrpZpVnH5iAM4J8LJq4tCyR3yUA
kr+4wqyiRFCUwJwMTGEG/zDBOrlJlzaJuVqYESVJrZO42sjiGI4iBzJNQbyTzj5bd09IBq3MayhF
LAJ98d1rRRJTNU0qKFrQ/R87RpAUv0ZmJHOy1jDhrUt84uc8l6cFNPlEwqn5CpIsLApmnM0LcR2q
UeGsd2f9cSyll4rS7SsBTC5lMWQE2a6jqcTu6KxbW1HmKdabLX3QvJT6YSwOrjIHwe7Ar18LhqOH
FTWNllXlhIopDHalXNprEPIRImCM+wXA+ew/CaalF0eWmNunoE9AY3D9/A4XRDZETW26DP2DpY8p
41UaOfX0UTcCl9neyawLv+6Bv/nE6fSoqs5A1g/WGfb5O6DdNZtmaEJr5m0rEH+sYf0S3oztppUU
NAshdvxOgAVa5gZ+X7/fZg0KMsssojEqd1qEVx3n1Rz5kilQ2UCettKZwIWSwShD5TzHdWb2027a
nEc76ii9OcjjUo0OWlPNGq4BIwnqLNONoAHI4Rtxk3se1SJhscpEcn/sXU4PqoLrSKlS8FpF2eSu
qtwDEdHn+RQNF5KmmGlybg3XZfloHhiWqYuN978fF3GWmID8TZ3lCWKC/DGbzOU1V059L/KRuABJ
RpABzMXvFQYQlqLszIUsiPIdrNcPNY9cMB9zaV0AUN5w7Z9JyhWRRvmRIiHvg5OOqk/dQ+hmyLLn
mLXk1jZcs5ZD0nCLU7LtYVSW4nDQP39j+ML77/KSAFerVDGLcZhew5d1cSRWtTbU4/lBBW2EoNxI
op/YK2A8c6PDmKZyCCO6LBP0iXysUXl2l3O0gcGYLXCBNtID8oQ4bnB+ql0R+f3K0No1hb7gI34l
0hTLLCuI4R8hDwV3068lo5VoqNCthzuvORO9t1uL5DiJQHqjY4jz3DcJPOM/mGBn4TeJc5lwWVwC
RpbDMMH+xy+UpfbRfJBcIM/HcFSbuIEixFZ34Ajljr4oDc1d2xGUIRTzbaldwvFna9aFhbJ7bZQW
8RcM9BVvqVXm/C4P7lfZe3RJ8U7JFIFFl4ei/52h5gSFREJiimH3JDcHubovCCjAwOIzDltK43yS
fEiB9OL/4F5gOuCrW0biKzmVDLOw97cRujDCokBhznovPcWbOFQ0gAkpvALIjtfq4ABcs+wzCr6P
LJzhOHbDS2va7En4EkSfcfYyMyyy5/eiUNwk4Pw5OZP6h+YMbjqFK9Aow3elsb+/fiBJ5vLrqiDO
VHVfvXsDhIsxrkUROLqh7DBL8R1qlW3EK5sg1YuLrTbw20V2weNNPUEsUSydIqAm2KhBO+rcZ4uh
I7IhtlPUduOaG9iX4nGOdrV98zHyF5/DidfUruBEGh+qyrv//LhAUDDTmPA+MafbusG37adYqe/W
+bx4q3MNVTeGeLfsco+wbDVDXFMTR9QhmvjDUvUDA/hX+c/+eWUvdEWKtqUTCpq3DDNPh00LMIra
4J6WbHijEoHJeWdSC7PoZOm8tcxLZB5eoJz3Q3V02VWe38b0t3Odzsc6dVxsYtZYyjzPNyeqdYjE
87eFOM0l2vKRnI2zLcC8ZdrAhmK62CyU3IllCGhpNFI8jOLA4+x3BYtVQ8OfsJSDksKG0E3usQqU
SdLdG3MS26EbrfJ5ix6iYLKGReWE9RDcONdb6mus8W2bBcNc/CA8r21lN5l1mZEZftvORaTGtPFC
Tmh53bGNsh/XICU/FEmXk5Dx7uBXu4Q2ruUpHxCSk1BU4td0PqWSVDuspWNyWOKnW5pHXIihoCOt
AS+PPiEFrbFEXZZy2xRH5s1BXqYO3Rb54ENrrVGbg3z66Guk5q1UhG7KpLvuzpAFgGloG6VeUx7Y
vrw0x1JuWn0mp4wDYpgciHHptU4EQcgqmTPRH2Ms7zs8FWwUPG26tVUem9y5PEAFFnYJNK9nVSpx
i5O6NIVwuvKZhCXfoJTCYyzus3bv9pwCuKUOxOi27p9ZZ1GrJSvwUJ1rolCkBMMExfPrURb8bXXS
GUxNMSc6EUx6ZoNSIxFHkucNez7c9V/+SLv67QV6Kc1lzHP7Zq9PDX0UsgOeB1I9E6uL6YJg29/J
KWXqnDs8UFRuU67voSrFBdgslcdANvgFUfqqFXQC++edjTYOxK45uHfOB3nlGz/b9+K1BrfB/i/l
+srTutJJjSSMOQbDFNc7iPELXdBwYqc6l085huKvPDyXo2BQlBq5E5XXS+Iu3P++gxI4H5C1dcHe
nHqobe3grErce5ZdyGwA80Juv3CdX3VK0IJ0pJuxry9apwODnXpKl874FM8wyhEua5AQBWNO2bze
PFHtg/bU7Xdz4ILkcdJrAvXC15E1VenkXgy/4LaFw4TEy1inxkf8v6vtYtgQ+7j72gVBGx6DpcRV
uvoL0EQtA97cc10SFPtTKvAaywATkUfLE0f6saeGtQa/oiFBJfK4yKQCWjivj3F5/+ILp8VvLN1v
dHpNJukgk7T8ApbtLDo1WsetemobWHy1tnm5oRMy1OHG/HVc9E8txrVld0bGkd0VJZUNyjIdo2u1
vgvaYzzWsuqeCmXlNO7Rxmy2VUkd11YVYJ1bNXRXS2HRma9GRivs0fE4r78QGxYnnpYhmNVQ5Iu2
FqamZC6P/DNGr4cm3kQQPiMLOBb82h6dJn8zwObU4kPrwOrw4DN4qACyccF5EoBb5VOtWJnF6aft
PzpDYGQNq2Z6P6XuMSpUG7o5ucTAHKmmqucAZmn4dR2Z9lqU736BOAay1zs6x129ROipsWK51Z/E
cuoe4Rj0+FWT1L6WFfT1fkS5d1Iv8GzKMnJg+NT/rnfnEu4zCXlUJWhfQbbtMCFv2UxCcWLCRVPq
lBPkr25V3Isq3of4EBz/ZJ8zbN//kJtPGBrZwpn0Bl0vH83twAntTccFxa03EI783ycWfHvter2v
ib4tnnUx5ZqVSS4MIJHmgVzF44xuUB72rEP2h23C3Q5iHOsYCfGYE6GynMUaljFkTrkVO9P0mQgv
zqfVKNc2u6KrGIJ4SIzjZtVNngUZbr5yEbYCB3ZglUyfTNf7/o5CK5tG9Qx4OIMY0reVlFjKbMvH
zdJ4KgMOP10tq7gmBC9ayo0q3O/WctAW030SEqfjL0A0MnTlQ2/p1QGr6Jd+9KnXEWjr883fRP5r
ktBRCAnujEgg/w3iikLL7AK5DtwsIXCx08yN5mZRh2yjt7O8MgCADlwOJmWw5Gi88j8TG8MwJ17V
iqN2jiXzDhZer9k2Hsq4CkAmygwER2EFOax0lwGGepbR3+p3DPyq+Z3cTdI8/GtGCSKAGhB0AHYK
PprecmbbSREUAqunkPedbqP0V0zvHB+N5cUv+ZFQJ5AEL9/7tEG4a09ItS2Cn79ghyahXWmR6nqh
Lxu1A95bpR39uUcCnOxOg5M4BV7/zCgsuFK1yNVKZuRSYc1YD0i3S2gtfrBNTMng9hOO+nrqHDeV
xAN7JdramGX4rDnM4H01FwUwPDEG83YobFiWIndunffS9ETLG3GhZ9LRZEXluTUbcZIvNvzsiTMY
fY8M9Nm8/nd6lCB5FmLSh2avD6XZl3gG7HIWDiCL2l174AofeSrWyztFVM8GJGQ2uQYQPD9FwdYz
+1CCszMVnNaUxKEEW6HdjI84qI9+J+G86oP1+Mhk3+5LmC7NjgA0XGu6TkM9NfURNx98ceDGXl+J
tp+Up0EKrfNxKKzB8BsNFV8+h395VIbqLGj1lwnyVnY6Pf03VaftBF87ZuaCwj8lm7SSKutk+RMc
xHs7GWd+gLh+w4mjrVDoBK+A0T83V91XhatOx0k2ttc3A9dMhhW10p7vgcZy3T6hBZZAonys9JjE
2ycLcMCTl9FGjKYAYua+RytWYcgh+uSit3D89MiNEqtNqr5iy4nEOJhEZuX3Z6hZLVpi5Yv5tmRp
XQKTFpM79WqFNkPAq1IvQhb0VAeAR9E+Nzm+1GS92OcSmOffcW+NwP7khVMsKREdVt9oR/8D9iGL
4L5P6k2hzrvhvRwxq3kZkzvc7MbB3wEXb/whtz/MeQ/R4dmF4XX/aOysb8DKC6sl8FM4N3dB+1Yc
ujbID0goekGphfhZBEurcMk75VDHkAhs5PCttssayyQwMec4ZlKGu7idBUP4TU8cXhwhLZuvB+V5
mOqucPGm1u0L3Q2G6c3vWLNmqAVX3iUkhJKtA9M8sxV0cssvWMhOvzm9rqbORF/meZC01mQ9nOij
M17G3zHbx1y5+3iw7+vtZkk9VOMwoWGSDjWA7GVSpNyYavkNXaGXJf19Ciniyp0r/0mCjM2hPvVQ
4ibxsXDQGT9BlxMlcx89uLWToa2vZWqoBtCGHUYpZM0ottcPpcgVPOQHW2HkZDnnYqvtKdk+NXdu
TUKFcfjlccJCIKsnwnrDNZpYFGggw8uvqlGkPDhwOoNOoVrjIwLeZqOgJBt5OiYu/IIEsbpZyAne
KFyKH7j7AaGqs+ZSFrRjYmeHsYWSoPMa5+eKKEnVyI2lxmPEnQNLL6yPELCCBHqWAxSCYce8r7OK
dA77wB1IXrw26o0Z97DtD9fDJT9pIGGAeItdXJ1J/dwVDNL7/YZDVs7hzHzNH89/Rcp8ABY4Nwiw
Peka1EXWdtpz1WHXrtCWM+2cTaIb4cy3GglOVHZOxwsFIU2pm1+ICho/+xiJOtEhFVvNpM2O9eSe
L6i6kWPaF4rctSpUzYUBv+yGjauuSAMqinvYiLeAc21BdRcXAMXoQ+bG1kLCDbE8qJKPTtX2KLW8
t0RLajneRh5Y+HtLK8oN2JGv4G9r5gfW2CUGoGrM2um9oqhjY36ABvEPno4PERJI/ZlyRvzy3S/P
aLnSz5PieqKXbzV/6QMNnTaQQdiIweDKyih0rWdSX5mf+43prKRBj0kbwqnWZxFVoiVKdwUQswwL
7j+EQ/Y+VMfjYm/1Jual24MROc7xzDVxEbVXrg/djmyX8QuhAoVgzhMzCXiCeHx2gxgM/yC3CoBV
/9tc11dMGzl3UU1RB2z9rx0IxhjRvCnKeMODy+8M0KToydw+9qpQw+vIbx5kvIWmzgjTWVa0cQuK
Yklv0kP4NfJY8oqNNXq3qduLyMHCdEW71zl4OP+ByMl4x5njLLXTsAJDbroQxbYeLBJ8bkBdp63n
++Mw/IvD9UHpfAHKcmJAn/1T6TnygyX38bEi94tJkhzU+4pyU4/bOv2UCN+O3Yrg933GvzyE01dB
yhMfgtYkmUkiQBzNDkSB1BwA6M/zJUUkjgdd5LifV/UhHmWS1HKqdDxTQYaron98O+y3rPx82/zv
Ti501xOxv3c1sSzLRBdOLACcRap6WbyrwOsdAFRCwd1rQ1AefB3l5liy1PWZhg3P73kT4C2SkWN2
cT69Inopvt3X5RM1bLMMMR2uGEke7jFjeyF4Nle+w4AixFKrV2J7o8cqB/zdarvtYwGVcCEInw95
fA5QThm1M5IAs7jSRFG4beyALcpDcpi0il2iuqyP9EylCu1eJieAtJA5jfrzPrTWeq9Z0m67WR5n
CAA3TQAXnTdauYFJIvjdcAxpRco0Ch/L4CE1I0TsE7REq8NkY+vMzZ5PiBwQ+t5TxleyC1XjLNpr
oX0evfSQoh/Ejsyv9VE9eTTO13oh4xAT5iYM4AbIcX2+ozt1gCtPZFucyZP8DVUqJrwmTVDAjDO8
Hb60wXertF69MDRmRDHl0iYK9kx6FQYCl+M9gm8ZdepxrdinAYROEttYfDgMNznqLFCRxCx7pty1
t+/1AtXnEImP84FsN6yDezhUf59yKxfLKOQ4hj9sXAhqe0+K0VXt7qQ3Q/uQYIGyFATPeazvkJcA
7r33Yo994lL8w5HvTIwHeUj7nLb8KDkIJJAVffoDsaY438lK4vHHKxMorwzrgIVy4hi6ip6SooOp
Lcyef9r6L43o3LZhCYsbJyrnqN8zxKPHcHdsFa6LBBnJYu3J+tYpZqK+hJg46+od7aXs6iANRrmR
/We9yaQlJO65+nMEvR4d0tGQXxuRvLQ33nMFyDvsNFeNTE3h4se3DlBz8V/cspBZAvtJWBfCkEGn
Kt026QF32RBIsZ6IP0gOe1N3qnH+3m5VEWNpqtaNBCZzS0ASaEWBKuGPsUhqEaIDH9jRbx9n5paG
V/lUoZFskFw6Ib/l7fZH9srIzI3Ii9j9/N1i1Pz3iTUbzlUNnyS87X8f8DCTuKsrBsjKZRLlYVFm
x3VQo0hJahSVXofSL3xeuVAf6pYVarEDVCzML8Yi7upKFPYPV/iild7LfdGZ1bEbxIpJ0y13834O
4JKLm9bmm6mEVNRQef5gEadxaKuNPI7P++K5O5OppjlWSlklRZDH6QKHbxRUe3Tk5zYwE4Lg0CpX
1RyvaM2jQVXpBkaaJsRyLofVw8K/fKKtqqTDIkeqfI2QIwB2rNBMsseuVOmJYEXnfuLpymcwTT4v
tOdbexSNbnQdrrc6aJK3FDvkRp2wolEHPnBdAUuR5U39hLPbzV6Mq5f3J8cJ7MIpAzLYUdWPDBeI
A4zMIQK4aFtAbTTUz0POmEgDo5zKiyre2+p2C8loFy5ZAcDnY1j9rTjT9kN0aegGxOotdiLR0f/N
iInN60bD+j90Cx6DHdHZ0O5sATZb44e9nA3QThikuNZEc6U8ZnM9sLYk/lkAIoXhFYHqhw9NG0W9
uynGSZlbJblG8b3jAIl8Xs3Nouyj0jbLD1pYq2ok93DGy+Xdhl/O1eYulWyCSsDnB7RQCip1FCcs
L+egcHZsKKig7jnr+DyaciBZit08S8jMa6/yHdOm3YQ+3xFU3I5SAz30sz4UJJarRV5B5TGiba2k
2Jhbx5RW+DPryHoujxPRHKecakjtaeJZu/lO2tXUiiFM8n9fRoRS6e8K94cibsuHA9UxKnu2DgMk
1kG2m0MbTF85/3fx41Q74XSNUVgGKK5q//xfqqA2GPuTY1BjPDpuUihyiopaQxixjlggvecTh2rH
TXLxNjWIBFYV5qtnRwHD4WHltyYzqA41/Mrq8RNpD1eHLU3bFAxbH9+8q+r8OwD1tqAtuwYVXHYD
I8srdYs8nwRxUvqa5JBnGqqhr/gOiBxN1l2Dzkm0sV2faHVypqp6PKQyUqHLJl5E0uIt+EUQN6H8
/TivwFZ1/ATp9s9Uog9JlDswWgunjWHfzuSHHVNeerfj/+rath4RnVbcnXeOEfGJmocDIichsCx7
n1G+c7aU/ZB0knYIaw2UiTRjf2ruiJWnhrcQ0eoxvT8af6D+O3CEHXP+nxJx8+/CpXmqIrVZtOqv
7YAU+aDKXiGM84eW/UqPTgsbIZ9SP7Rom0cdIkI60UWwdkdX54eIXEBjyM+bjL5oPm6ncj4cOLLW
QZHjs55M8tEjG8aAulrY6Dr07KcLZo6gVbn9ffWDYnXxFd9MRvglYI63LLPd28vIWGTTQE6RjEUm
fpYIWnbL1lkiqcVKfL2h92Jto1Yg3P+oPiCbBa+IodbxFjPRuZzcI0EuA4IFWfNS38Kr5dHBwDQx
TpdLWewWKj27KIJwKS6i5+D2fMNmE5D7dd9b+heYJZ8uXYSObZCyg/EFNIxexkQEsuUEoCkBWX2c
GtUBOjASLGx1jgk41fitBY4JXVKfAYnPH+w9hrk62MeFG+Nr1XrZ9C4I6hqu5djZKEqQi/+3+s58
XJcTVeeqMSdI773gu45ufj+2wqZo29NHkXoBr3T9VIENzHdVfC4xlxVD2cpc7eSp9Sq5uNJsx3xQ
MP1tvJi9gAWnswU3JrQwfMK9mZTU6tj14q2x+ZzYKYp/GJBdDn/04JG75NqkoiYWBOWkbWHNRsd1
sSzo+WE1LHt/5BlGRKvOvv7PV6wGRTWzdye42Ck6EVHIlESr7hKSbRoE0wYkrSUq+miluDOq0L9P
kVe31u4+F5IMV2PIY8iML4ZKbNQSYZEFJ2exp9DBNM5DlLlrzjOyAioL1zdcTNraeqMyY+SVoEKg
xA+C2qJhp2Tk4yVtHLAUjnC8mSf2CI1ZWEfv+WZwvqfT65UBpGWIWg6MkVi45OJdps8SOVEG/wGD
1xvWkgt+I7sT8Nq1prcSNes7L5tu+AmZPfWWWPAssTfPzXLYbXMiyH7++6H8iEDB0uAJsjy64VGh
/lTxTV00oRjsv/gz09nahi5YxDJ3oXM/dPCjBPcPcY7voVBuRX/ydNGEwEMGCNqH07aMGKbgO4Qg
sJxwdaf/5Bp7zwbO3MmEsazRe2w1sdVfdb/g9ZCBQ2U0lC4wac8v2P52UfAA3hxxD3Aa1Bsm/JCz
hJhrzZtUDj9gSk3XWqecJYcR3iyZGEpybJQsHS8qDEtgR4LP4c5z3AZXFV0DBHV7C0mWAusBSpFf
UxVGmS8thytmOtRXOyvz3r4ZZe6Z7dLpidTGvxGbiNJiI70M85/uMK7jmMbQWvboQI84jl1LGE3g
fEqf5OD/Vkho53VAV4Em4m+ng1U7vJco0h9bqokSTM1HoGgMkh3dLk6gFxK8mYzFpzDr5eUNfEKV
wsjDo7dGc3Ux/YcdYC2fgmjeQsx6hBPnEO/dZiOszm07qbNB/EnGW1cfxjCldBBcCQRLBfeVx6Rk
mCJQ8CL62EnQMooKqb2CR9atLndwEToQmuv5iCiY1vH7GauCrFZHumhWjp9N2GI4jMxFseNqU7mt
LzDqw9gQ8dUylF9R3N7bDmitw6NNYpBZTB2MR4nD0kRnY591dvA7Rncx8RlZM+oVIztrubIJ9mG/
CylBS+ucmUaHGuzhVG49b94VMFpLJxAhJGBUacgjjH04OxUNSI2twdJiby/6EZOmmtYkS1ZnQnTz
67iYU3jCKwdPqYTapWhAgW7q8A7C7heHOgjyHXAUU2Cy/G+9DSy9PvwxUijHIrYu721p8pU/hruM
flavVydbdmEXeJLWm9Y0uMVNB79OrPuuWktqLZr5993X0ykaWmKl+vAea1EDUt26R+zdPgqhIm1e
BwKqY9/Q69+Ni+6sh7sLoKnzEOo3Sa6eyR4F/6yJ/O2eltmew+M84ApOrBck2aqg20Fc7cBTzXwB
zqtBMUIRK+3TPHsLb+e319eRqZ/eFDVjjCpmaSDGhcxulpJOkxvF6H6NXXElxFa5fU1HYdAJmuIP
HEQQrhbohMmfWEuD6ZsHPcr6uCLDKV6kPu3InE8uiPLf5gjw5F0FOXNPGcIHYTLSEB8vpY4BidbO
PodWhLDdxWlg2chV81Ie7th/vs4PA8yIcoy7rJSNnqrbmL3iYgQlOnFdxsoStit2HcbZDX508IcJ
3FJfO3dabQgdK+aknji6lk43ysa4BLFj8NyUCtwGHtEXCYtXl5xHSyESnDrYfOkBo5m/28nQCQAD
/BTDfAf5XiZLcz4LeLQctoM6NfuR4HQ+Vg3cx+RALp4Q7JwnmGgrEpzmTTT2j3k3wI0hpLkymlZM
6/6jylXC8jVsH+qJIetKAGFSX1BOCBVqwI7psOfXZPjIlfNLX4CmD7pGOCL7aB2Ra2t4MnIUirLm
ZWj4n2/B5yOwkzVPWfAxmRlLdiyaRrSwY745NiM2vrpvuBrEhNHDh3Rm46YjVbYf+UFv+foltAuM
mh2rehTnX0GLQ3dzveISLsfsCnN1RYoO8oHkYT1x1PrYlX6+dspAK9r02Vl2pZPb7IXUg5I424Px
qRGTvUNfOXD5j7hHgdXV4Ecv3beHL6i2mX4463Iv7UJp2V5KiI+DpC84kN4sVLWz8qkzZJ+nGzaR
nFgpIBDI5d2KcxVEYjoNCUMyoAhZ4BrBPDirS71dyOCqi/tKR53nNSM9xR+f5IrHIv1IU1a+ZlvC
/zqh4QRaiurStIJqX2ATk05RxInf7dETxiHWpR2Bn7WJaYWmtXUs4T39UPlefi9P6EFNzTdpYv5u
J+ce6RcgM49Om6MCBi94l+c8lZeCqzaHD2iPhZfkcuOoYLFlRxX9KnelqmFIUxrKwaPgvgDeVtHd
p+nnb48Mu3cR4rzogwxsnQ60YURSKKUdBV88goHiYlZq5tjYit0IQbs5Lnionlxt0sW2ctcndkLS
SS0cM2SrFzSHUNMecz6Se0LUr0piG9zCCw7dqt/iJGnDIQCYr/S+DRDDpSe69YNTDQNK3eABKUM4
A2cMI8uRddaVcBs5wOq3J8HavlGHvwPFFIMuemZqEJR+2b87k2oJoxLGaoGegn5eIC2M+osWVE5R
Zp7F2WVxeZSNBfsOx70tSLPSAucgFvsprISlniUsQ+sFppm7U6wDuFNO1e584fL5IVOKU/NdkkWn
Z0bcFSwM/wC+mn+V3z2DevoTtZslr12SU+fqM1JrhvfJ634fzx3Q5OVKUNPk70CzNT8oLQd11hah
5TwllaNaGeKCtu9+6dRDqO9oDgeKQLDvVNxei8D1Tt0dhh+QQzhhIJoc/X3f0Hr8nT474TCcU0i6
BeU7PZswG/UcoJ82A0Y1lN7lHFeqcxv5mWfpXp2zX7/8eNDOyza0QJA8hH5gpGa0k5lTg2SGSpCA
Y42qB6BKv02gBetpK7HD8yHju6aEvElzyE7ulAH9DmFlmrxaGBbVT0tBIfXhvd6t7qQo8zPHbUeZ
5yOZnoS0hNsCsjYZx2BuNyFz04EP2JlVqJdBYrrk+zVmsVHhgMoDF+04DSYK+UNg5vrt7EGCeDFO
jGy9gIrKLU6C3WOW6LC0JQqWz3r2U0Amm2hLVbz0LTMhErqcdMbe0FgAjJOKpU75IXy7zOSaf59K
Tyo8uPJ/dTQOBlHyxJLFiTcQ92ABDQWxc9Er/t2L9uuYpQ3TxHrpW1x8CKdhzv681rKaZOWuNGS9
/pkUbsFo6/g/QTxMpJ6gG1lZffz0LDBcTHvZ1RW1sd/1/tQptA1B1dHtfSuur89AsYcka4TQ6yOS
Ebhqc5JgjjqCed9YomJvMtCObRnpJcz9w7GDG+HClkLGq+JMsyjgq5CB0i8qjx+LnPA6EBDFBwd+
FP3w5BfCdT1Ct9RvFL5so/xJ+4BlWwIDazCUBH5NHBBu5wqSUjOyWP9Ma1OfF6Yz153+7IhXMUbr
8qRGa1PAPCY2bnbrE0+kYFLFF7PLtAHN5MCRhvrkoxCMql1eyAnPjAMMbFGtrgXdVumQ81qqZxj0
aWCsgGKwmtqRhCFHI5ZerauEULYTJI1xqSzgyflqWS/MmFpLxgRT9ZzgU6iRTAFwsLpTZ7GisbNg
ogaWHyCgbpgiWDE4AFhpctcRE731X8qj7fJMIFEDn5WeOXBaXtmL6B/l95HyKO3XOq0mZl3/Ta+1
SyoQEx8OBYgTI6Z65oYrTxR7ibhY79964Cxloh8MqR2lnLK0rJqKzIhkTLcLEnpGXU/WOhZBD9wQ
mQqqiylPxouo5caFvUxQfjMcsAEpog7cX0Lzo7HpZWrwlFQRp1LmpbClBFPRqgjex2mLHFg/wh+4
1eVL3dpCtvrbRhNqcK8PdeiORsvAbLZhED9KTJkjkvAdVq7ZdThlHAR6u7ZDGHZ1tCo4ZOnDT9LF
dnIxUBGEI0+rN6TMSrRDaCh5iYBQAdi1d8/6jjg20GmrfBvOwfS/y5hqG8bKKz/oCnIOfxRqMOTt
exJhomFwyqDnTiv77plhRZ7Bnd3S2rD/xNnb1YPnY0tyRY7Y8ZQsmgzySr/IQMydGlPyc0TWc72g
Bc/bGtQzc3WlXgymKCGFDGy6FHBVDP4VNN815prQyjh48IDT/Oc6764p9NUo8ErzBNtXxU33mEZ0
qBPQsO3dIwgVRBBqWbtBIkbAW0nA+e3Wgm1yjxy/Of5Rf1S43oNgpMyEXn2sQabVLYegNv7LF0wZ
5wl1CsiHtJwrNxtNe77ZjcJJbNVobdbPKLW1BpLApPrOLXgswvVR0RPWadXls8gip64W3EqGEgsX
6Eysdj9LvL7h3uehZdpsdJFZhqiODWL2D6d3jYLjW3znLiFQ3ZQ4LfWxYZAZumqr5goKjoLDNHQo
C0Ef8E4VSik0LOQ7lQEyTf7K8Ms3gHGA7FJvWt8FNrfvDceiZ594vL4wm+7h1Mbbrb6U9b97ODGL
o8AbRTavqmvO+l3FH6l+kfpFte0NQU5K03OCH5lmTVFfy6Hl/o3Cvb6MwOl6uEeE4zNNIO9MXjLX
tmEwI4wyk/9TiRxov1kKGGV8yqQy8d5Mk84HMpDQj0JNwmd6QF7uUVDGImXhrNQ2n8nuzdeG+9UG
b2fewxyI38Ke4iURwAOVvsVZRG8yBbUZDmHqIHpZl/GqnOjyJnPDWnKAgwtt0cb7PYfMcTUiN8Eo
iEiR0zysPOkqsMI6YYubWECyGKL1dYOjks5nNoK3jeuKwzHxazFuKAI7RJditDBb6fKppTpB4sru
vd5qUUHKPgm4Cs0kisUUjCwb91r/cpoLWtUu9hllaaT6nlQd94VrB3bTVmXUJcXtiPxIJJldpKtx
s7gdFLoiRH1zVqd20uPorBD0pb8dDAEkICIjTJu0e1NUKV1Mnwc74kgvNH2abKZV/fd2sBxAU4EV
PpZEUMjUTFeU7if1+DwnpulYLW7xBGFjRHN2cWd2gzLuD/iKnQM4dShLorv5Fzn4x3CPcBwgBWXY
uLpA/e4/mETAFA7sSzm8jD6xp1JP5G/Z9cM3XcYaajjfMLNYoSOVZ/OOgGtXQL203LuT/fKWKW2T
wDc2gpQmbZvdKPqQEH8BYw0VxpjrfvXALhSbsZtZAIrLsJuy4pPnGDFCbln4s0RCo6+uaQNVhVHW
iYY0JDftf7Uy9xAQ3Yf2CLbnTZO2P1ehXgcInAMOhBORBI1bzNn44uipTaTczQ3yA7Z07Mst6x5T
RUhCxbdT9mJjBSv6wt8rEI3I+WnnfFshYeOWaOvO6QXyDoPaetAZUgdFWqqJQngVL+1/BVzJms5W
GmyJ39+k6L/h5IhGNgR2stpL5E8+bQmGjBcq2E0DIdFoGBvwJongaTSOcYZtyY/2wGwutdsWk0lX
85kxnOFSeSzd38Y7QZOwU1QAbVTkTeosrDs1c5Qb/b4CGBbMxD/AJf8OI8FM6MKVM3vZ/0J2W76Z
ShvPSLUBk41NUFupibud8CaNMRMp1C2DYlkvUTtJpOKJNlQG2lbsao94YjupWaNCtW3tgrtKfhhx
taPRDaNSDtEAVXn44v1b3PTBRCzpj5Tezw+hX3QkZKCCyCcfPu43fNpzggZYJqYfrosrg681VjfJ
iD8VtIWNNdcTybcXMBDY5T8FsGiqbdM/XLHXE8RYTaevSGxbbfd3iNFWDwTX4qzG8EYlOiYQpXwu
hDXn1k/jBpH0bpONhCebFL3l/CdDTVarsXt0KPWkzH59DYeQffUo+RxUi0DCkTx+3w5RQYWLA8OE
j9YHdyqvMHbEZylEgrlHiKQmNJnxQKBd0wEuHh9vUcns/ZdpmCvQhoZKnIvkb1iUDBe36IRupIxv
AXjBe6BLRorpkqv48S3VylffzsGDuVkHftkVWetGIjURF4TSVhfPT28cYLKmE6X85RLA2TnsPcZy
GSMFAmO6QAi5et9slcS8u6fC1g4X9l13qtlG0ZRrYF0yC/k03xebPalQSTHiBL57Av2vUttCfbfF
0e9n/GqnXJVt8EMglkrQn5YQBltltm/0iBgnnFQMB/YHuWwcWROLX6hu2/l3iqtD8exd/AqVPM3S
NqHWzGFDED/1JRhjBP9y6EGoB0vwjR6aBRMbGGU9eBTND/Yzc+yUlMKplvMd+v4NjOTUNmE90lRV
gfWDVU3F/VOvEWPbmmInYr7ZTl2jaD3p6hqEX2EnG84Xzs32ctHo6+5hqcSl2OihcHbSbNEicu84
shWTO63341eTo2D2BT8tw1DSIj3EnZQR0PlUlCWX9Y4yLslttjbbSyxzXz4YLHShI9l34uB4pmmc
9QFt3+LR5O0eebr40/qJklQQN1WLy8agp4UUGJUSCC0MOd1dM/JzdyVcgeeevxhBGohju7ASxkbd
KLyCbQGEvVLJyFMZcInIng4jESYu6zxxVMDaUI3oSlXmxZA6KfbgZ1Lb7SyPWgp2mB2APd0g+x5u
GQDS8egpXxfJet5H1TzRDU8tpXAhjZIBtjsxHgknb8EWnSDW7fYbMjS8akY+eiSpRMoTWcrLhjUF
ySs9tflzzyXg1zlDjJAesRdIAcWXCOjiYY5QtgiB32LtkS4kBADSlgMYmCDijmlUjAqWke3tzeRB
A4HAxWFpiD2VAvGjoEHGbCpQ69vxH8HH8cYrnQ9W9mDU0hcxEhNL8jTtBx159hcDF0N6itX5oa4Z
zu/Tzo6TQVo89epdhows3UWkTI6AaOhwiIP9Xsa2JosKwS4i9yW+B/xXrwLpaPPmDb81BHroq+nc
RPitxjZEhy87yO1AwIBcxKWmqPSUXkmU9W2HI1b6guTOMtC6HMhO6/zXPUYI8jWUbIhtWfUxoqiA
/jiobfKbT9e26FuYGqSqbxrRCmLPkZLY7UN3UDskjq8YXBFjjVg7F60kMgsojqEpuY6Fdl3sUa0O
IORX+7j/oqqZUnPpFDYgCk67SLKQPTng3oADm+/hY/+VPntXI/lO6ceF1rC2qU+qA7dxf0L+9Git
8Axm32QjrQ0USN9s5DYbTMCJfzzClw2unCETlfbDqNtuH+pv3YHgxXdV+pIoEWhS28H5fgWabZ3q
k9rByOCAeP9mk8+ZZ1Hk1WhHXkd1GSm0jjEOATdMerBpQn5393Ir+M+yyGn3BxIudFootkQ9R7Zx
9Y5BqBnbBrx4vPhcrqtf1GB2Nn4rknlQR+2jO3vw/ZRiGv0zQs1TdXeehDHZXYMreA62LXbb1Dov
fvlBnPYwCV6gO2gEfCo1FK/d/FDKbZsU6YflQF200GzDZUB21puZHiulgObaJsN5SZZahP5j1bU/
/6rbVsl0Zx7nLbTES5huMIM05BrJ0DimYpTZU6veh9m5F6D2lx4Y+MAi0LrOH6ykCcwT46TLxxHB
JfMxmwTsWE/VHlqW9UZD/Lg9Sc8Iqy/Py5ah8WkYiXJb1WwrYNe+vcX2WaH9R9NkJlkTqwnc0pYW
Lsf5xwcmpOMJ8exkeyzH2b0xCgntNqcWy/TJmIQQr+6wpcJNEkIHmUHTviBp3eZt2jKSnPz0hon0
2gbHC1h9g0Brr7VEwTWyCRFV3nT6gadMOHCuhYdAePHCiKyZhHyNdqR1V/o8hb+NgytpGjyI1MJM
qVYshbg8pRkgib2lt2UkvQhEm7sPI4ZovWYqxn3vIAMIMhVksflNswkUGTDNqlMwJvLmgeqGyNJ7
a7x9VW1R6H34eTsWvjyYP4svp5ZEZN5glzS1GwkKpyB/yInI4xPBcct3QgfQR55jMkm230t0xaOg
rsQm7xhQ1puLYuyOyVVgjcLLc3wPrHB2iXAbA4XES196o+whpl/tE8DU6PnwmESFd2f8UvGv2AJa
8RQddMRie7a1A9bSDMMsAkS7dlVEYMAdczB/WIgKNZ24glWP7NKImgBTg0M5zjVIVjaIHUVzeP3e
6vNrqHC8GqhRTEf84sCoPLg7OOimncpYocXc1PZxsu7CU+UclFXuhqU4CD1z6BGiOj6iJbq3/XMy
WF4ikWtHIb4U+/W2GWvI9zKJBehHQV8JyX36645kYUGIlAaFbjtlfLdR5XoY1MopLLg1RGt2NA2O
aegCLe6hef61Sv+P/z4/lp56wNzdWY1DI/Xp159SF+jjJnXJ4Q03mT1UiaTAUKwS87N3gOeXUWkE
9g0mfA3fOQm8WCaZ/4hUI04ZO/xmb7TFpb2TakwbadlJOVxqRpFWWeiUOnuAB/RvmPf/OHsXFq8y
5CKx9zJ5SV9/JexV2tJLSFw8XWvADyoQ3zs++KqMztM+wF+qwbUT3mXgjmtc6LRe4abS28g30xsq
051u6sbQ5j2Go5IoASCfDuNVrX6m8shJVwVLk0zWH/iGe4ENgM7QcPmvhPEZBiDqhB1MYql5aswK
0Ac2FWFQu/p8UwDU/aHyQOTgHntJ0oHV4eiaKQZbWmql+R/1tNPXnIdZMQyXpS3g/gnLRbgP3qDI
RMqNM/3r8A7Ie2C19kjDvt4bXGIwzMnp+oJiqwBzPYqA896r2YQD4tcqxNUoIamIbFLc4UcqH4TR
PfoPvqLncBSUhhedPi1zAVocNBsiLcCbKCt7BJgFZXTj8if6zpfHHA2xVX4XYU/FTWloTfmJovio
uwTxTezi3JwqgSDevLnhIxxdmMl/rdijEoFnRe2hcdTWYrqyfK6q3JuhOvqqsJKXHUM6TKAFBT0n
2Ta1yQqVjNKC6Own8bw6vP7DV8u4uhccYg+XdX687yvnrddqyrVfO4FeAtaFtC8wg7ILzUoPd0AB
5YyUPqbK5S/71Svuht4DiMvvm9UzAfdVTXtLNS77L8H9DuFqFBBB4tHBF2Y/KHk3sxrL1+MLBvKB
75WCXZWSEiZu44cazX5HPfKDNNnagx6CXDVKglwOvedHuCLSjpTAPKk2Ka5vWib0sudLDB1apmrn
QKiq8EkfZif2nKVAWjqSrdBiguZh4opetH7XCen5SSVgXj+2BbhIG/EJBH2LuAOQ5CKscSTXClek
6XVl10YRicTccTzbp5JvU79atzb7fGFZUeZHadSF9oqjVE8vd/xdS1D8Dl0/zssNOTSmDQIkv3sR
9zk2rpEquzetPLwgnMd71zbWi9oMPd4MMTJq9J4i3KgnJNCxOVjh0j3IL7pKHVK9CjINxnvDuagv
xPsh7O97A6+gD1ihql1HbByV6iYCM7SS+NnJIGWOKdzXT9KSMxb+igLlCWxeB/CAWP/dbGxScod5
EAGqXvwwb86Ox6Cyx+G6qUXfIuziGlMu13N9TuQXuuhD9+wTijHhUIX9TXATcWt05eRlKy53yYRa
K7S10KVjfMhFSUlsvWpOAvzGMUEbpcQhgs6Ox4d8OpT3Ser37H1IRGRa8UI2neU9HB5us2NAHZi2
w5mDNTnKvkp3VO1tK/eeNNUzQ4bT8mI8pS1f2kXoiM33q3MijpwxZEG4s63BgFTyVwld7g6kSdwf
JBp6XUhrWRacLxS0dvvlreZNl4lZ3jyCzyc9MJjuFYoBENVZh6wlJvr5vvi5dwXduVw37shEHxbF
X6n3uzxAjrdBZzo9X9vEJieQlJsVXJSgYneZ6mC1bVCCNXdASsZdl+lQN3i7Zt17VyZEC+5VxH0I
v17+EMNbK2yFj2+GN1h4Q67r3jkm4eHmV9nkI4E2b3fc+iwYayPWW6oyVfN2Rnu8JTF/ttJFEn1p
5pecaz/V7AllI6N078vuGDgXvkz+jZXC9Lvnj00wdFHWSTp1t0Xl6Wz2cs9Err+raVRdoC/Jyr5o
Xd969RuoX3D93rJ+57zf1fBrXWvYxLfMNBkVEcq7szUkR+G0LxH0Ns9cesscyJlQZwG12KIQcgDu
k4bA0MXpDZ6dal3TAlkWu1BNijU2V5v8lQJYhLwID44f4mjPPNJ7CiLWl6yjIt1K63ZSFWKER3F2
zMTj31MfDfUPGHjrlO3GeaPyrGuFv/G4pm31cnNgj4cdGh3jMGTuyBdnz3FbMTxhhzCYOzhUE469
4pEAKkkn5MEFhkc3Y+3s6zXTQp/pAQZ9fpTi/yHWbBpT1JQJYaXM3HlXl5N2Sa8cdCtReaLWhVBf
3961A7Dmoo8WfmHJx23tnPK5Yhp3DZIn06wI1Sq6LGckpnnTKO5jTAJK9kogyynSJVRi0JGypIf0
yCFSkK3XlZF5kzQ6XBeMgyZREK+HDDFvNWhu1ck6CTt+FKxYip2qZF09+zcus5dX8VzGAJ9V3jaw
ZB9DEL1Ih4mj1bPg+m4cQ0mQRxB/2zZ6wwhxARbHVwgks7/wKskGobqj7tUBWFt3raeHKq/5rqoR
g95GwTmAofuyet9RJaldnR5k4D1BloVyZa4zkNGK4VTMG98dtaywUI5IZAH7G7Kon+CTJi/0GcXY
8vIRP2r/BLOSqnh2V6Ms9o4VNIVHe3CfanFxrlS7v1LVI2XlTEu9PAM8E1IUNAmFu5FmbgYspFJ1
kmCy9tVTM22/nXAmDaUuhJCip6Y6g2IxUcdezi3H/SDsLitVo8QPcLuciegeJfZk+1cIJhF21zbP
XGrqQwgunRv6UGG3qmmoo2yjEWgXnCwPVDXh9hgEv/SHGnknkglvMw9Nfa5Co3tv3odJtvAzzF/E
1uBp4OXE4MsrM+6tKvyoinvYp/GZDjyrecyVnRO9vK0lRm4SZRuwqIyHlkGAOt3g5nDRrYZrlP2b
biJcnDsPJ/i2FMvCsrfjymfog7OuGttsVZoboCNqG+VXLaS78Qb0DC3773Y4jM+pM+uZnmCf1R82
XJefjOT8iqu5jknLGwj9G5CCO7Xv+Q5DoNfYwjcgsQRr97hnGCxux46Hx+Kuy94cxl2Oe4EcTk2R
QWsnJu6VeXTuSALk/Iz9Lr24Sr8w6rF1ppckk0F3fHWVfqlJMwFPvP2DE1Vn1yyjRK+tTCstbLj6
r1vD/5dKL/Qju6AD8OPxEthzZMBzKyLNO6/KyVZA/sTIHFnnPEy3fz1BHSd3YLt9y9iOfySwii43
8uF0OlbRTFeV0fk/Z3N1DBXOoPAMQWj48W4rWqX0HIO88HhQ3RETxMrWYY0ftbIWKI0oPHYPXwBT
haWtgkLFjbDgmJopk24BXf9R/UQryuS4ohmdnkIr8zCY+Sbq5Kg+RgqhzyjXD2xqp5hQ0HKqxNzU
eWFOmOxbNu4AlBm6WdZTR3uxg0RkuJUUKj8bPSvFBiXzJgGHa8OmqeN+ENUA/cr8Xnr+pBdq2jf3
2hVKZk+EGqmcUC28frYGJ3EJG8hqzOGyVqGufGRo4XVAirJ1R7w9aEiN3v7D8iE7engJVegzVK2l
+R5B7X1lea9HxxGKOKXHOzn5jG+6lWJkBVw3qrv4RF5RtYV2uUOOUm1Zao6vsyTG9VvoRE58Dxa2
S0lQwvQuMnMMybReKT6IY2kysJVky1oqFweS+G7JA21MUOzRaIbzR2D3RGujVWmZkddlMq8FiNDb
oaZJP4O+trJaywRfLgO7OS2hz794r0uSxA964mG2n6r+pRm/wG88sVpN1v3UrxmRO5JIqkr27BES
0Ey0YuB3yoY3N8xbIyqlm0c1JWf/78A8R7/3kwVRlVZJWgLXHYW5vw4ZLIrVI9VHPGMkDH5GlhvS
Erfvj1dcaqTLDzmyV9PDKEQrXkrQ2mz9n1lpTzSrWeYyINlMwNu4ijO5iBNwc8zLlPfDiJIoK9dh
l+nY9dowp1jCwI96FujzdG7jCUcl8lYSpO0jn/RhLuzFCNyZHb2+KB3X6w2mxB8/fUizsYL3iXua
4pym7p9l7l9msH21CwzriDoIScjvIV6W4F+SJHWWN8CpJftLJdf9o98yDDhxDtLBl8E/OB+ntyPa
wSzN/YqJVIvdC6xxP+US22Vp7146/6IpH/UoGglrkxOveoPjn9XUP2zas6Zk+PcfU0G2IicjAvKo
pjdSdOZxK/qPHiz3ddgGs8l4TvlyRnKZH6V1VIsE6+aWBNs64SPfcH+6V0lOTpLG+tN2ZsdFOn3A
o7NHgAWWneUCtYMcZ0OlbPGbifogUG1ARix51/2BaR7C/3VDkQaCb+1xAxlIV5gqtAGRJCmgAos0
4mP4yrqr0CSKXcHV50UZPPtAkmtsvuj8Rs6XtZhzDErqYKCne1L/RBrGseHFs2dgkJPhXLFbKJpw
q24ayF0NL3R29UV6FEo8+VLP5Iuebs1EoyVIn2t1ywvoQCqXwZGtKxC9Vsz7ARJ8vuvrg3HCgs+R
zr0IfshS+XcwJLqNXob+BT503VqUDtMFlqCPhJhnlq+mm3jjqvGJpIU039HpCCtNK+SjLd0NhyUN
JnFLyz7i5Ut87M8FnCwpRtfyi6POd9YZfA0HwxOII6G8tZ1kYrJVhCGpPEPNU0HGUXVMfGYG+bXh
htEuoDwV6Flum0LftxvxsBAqMlNnfHjADoGdiZVWLXTsEdVbJeUE9kd+bvN97j7eQRLSkPsW118/
l85XkcdaOxCxPua24q5tby2NCAh6YW3qCF3vhYtIaeBPBwcKRidGFHdn3mBu/z/keNMOIxiweN4z
Ln3e5vfPBXYBlFfoyUEM+VSxGMM3O2R6NokVx98c5qnI9PDC+9uPK/oOxvFEz38iLXljhwxmdJES
s/RZJSySA6W4QD+o1+6lmakUnO6fwEy6/nyalzno54tgF8dDugfqZcFn1KdGKjduTfF/2DdWPTsl
XY4/B57R9nW1vS7aKvaACqnpaHUN3fH02iAsGZ4Nt/NCcFyIsenRUXhB3PleqNJr+FW+yoAJbyQs
ItUp8nWWA//M090ueeQHZjbvZeUr0g5Pr3U2/Uvn8i3U728auOLOvdu8EOCd2BMuwsP6Wp0bMh+Z
gwYK/NuEHJseiWv+H8cLshs8T6xp7tlwJNUzJUoYOtWVUUjXT12GMar2ZknJ7b0IbKrXcCD8xvVX
7aUbeRyCQUmL6GXXfWHhAAq/GntKpXJn4KtPoxz5Xwmc3uhB0077dlwe5l5Y+fingxMCcoZ9i2KS
seqD1L5bkOzV3JK91DiYodQylH7XVHXEMWbW3rUoe8CEUft5aMPG06tfqDdf/an5vg8/eobr/NMc
XpiyLwldphET+Y4y0UevwPJAHmoTxGIv+Dtav2d4W5F1drhhf6lumdVw5RbY4YhX+NOLTE7MNk1G
F/9dI06PkTTeYUgJIBAjQvsiMPIJJOvRBxsgkTSRLcIHsL2kjWajqh/yobWPGES188K99DDLA/oY
MRilOVnGdk7ngm9Mw30cvs7Fc+1k1VlVzzo+t4+DJ0Tv9LUn2lfoKyjEPXttAysstPwIkz+R9nFg
FfT6kefU7VHrNvFCPWflt1Dnp91AxXsFXIm32kmdys1cFoRvJcRsMepoW/fR91qsP5KO8ocVu7Q1
/cW21RS8lWmnEiMtl2UIUbtxy/ZpZGIdhZyqescMKoYqaAH4pXJfqkAqi7L6wrd9sZbuVLxj7Jw4
/6frpSAsmOv4ATT3va1kYYkpnS/SkdMSImZpMg3HTEK9Ap8pirOnNZuRDz0rG4wa0UXyaH55i3iC
pEODwkLVCwgMPN0YIXjUd/kzFSYy1cmlQJj0Pp45+bft7rKdM79yhboMr8eUK7cjWYMStokNa2LE
n9aoYaMuV5M2IJCT2aWG8OwvrDhU4pFRKcH8JsrJc7T5kFZ2caOPtibJt8zYfuv+JV6OqbpaYcp5
Wf9/Dfmqz0vft/00/NeFsDO+m4uE7gdaaZ6RIOupwtW2q/4uxKngXGy/1NiMx+rGW+XIfd27L0zV
lH++0xQiintKzOqndWjyHB4Niez8aH2jnb4A8cEVs4fApsfq1u1nI0cS6vKEYjMtobXgVshGQ6Bu
2Q9tluKpYiyfgK5XYTJQ8flJLJzq5NyzBVqcdMmiIR9QMo3ag9UaPodTNEiZ3VdDapSKNm6Y0fKm
zins+5hZu5YdcXgGOTMJIj25EzpgyG+8FUW/uqIr9J9zI5vXXLFOQBdJbNKn/JfF3RDd5aEYmFLZ
61w8Cb/jzg61oXvwharQenTApF1f+6FZXEeW6c1vosT/tmxQ+0gP/Azm3ojBAzVeEgCrYNZq48Rv
r82QA2+HLy9FDnEbsG65gwFtuuiwXZNax+KT0UE7P1Ls/boZQb8ypZQ3FYqQSD/XEO3pSyYgR/gx
dwo2eCY2WU8tbtgrtaLfR2q39dQT9jsAKK8Z3DJIMVhn8Ze0YmVMfMGsZWfbmkdj2zXRWaMH7RK8
RDAgk7YQ5DteFI8pQdv7ldXSI9r5SWuhA5/b/bPwxwH+hHFNZ+XARsRZiXZbxicCpN4viBtMDyYw
fHcGgSCVyoP/gQ+O6PakUcDyHMV51OlnnYpJGJIDNj5WXRYDWN9aTplI4zZ8YfixHV1W9iMxth4B
Ohm6zsj6+yhshBqaQ4v8TwbkBiGxNuDkpUmIMq/27szei/w1wqEpcWLnjCHoKn7uAQW7pO5sdjbh
kQtO+hXpLwXgDvZNCvNSIutGVjKOL3Rm8ZoUOjxnTed48+3xiS3pGpkuxLHjUyfh1SjJ4axIOTPp
JtgLddQsXtBdfLOHlMi4ZDIv9yXwHrEvfXvmCmS0ZN3S3SGBwovH2PSFZ2+Y9GZc76Aa1Gk7AGdy
qc8e4OXlJubViVkyxdC3PjPZ0kn97tH9fVGNvA3K2nBB3p4fPJHGHl88CbcO00y/Dty+QKobuyMF
mxXN2zZclcRJB7NdK9SC53E1kQ4sh5SLnfkcTYDBw8ZJXyn73FeI/did/EKzep0cOGqeiLJdgRo1
VPnsKGORUDt5KWtxjml9h9h9FyOmMNbcjQixQVWGVFWCxGXTH5D2nsncfzMe9xiPuOD2Rnscemun
c39mcyGmMEpKy424KYnID1poitQyuLA4rZ2COckiGL9TBUvfiHSYTwaFW56/LMJm6+PzL/L3BoAQ
7HNZnnsdanqX1Tk9T2HK19B8f3KDA4D9NzPBChf++dazEb+ftGh6yfXxSAeYbZgQqbDIiohikBA7
Z1OEbVTrjCu2xGjn2yxUkxuUib4piCajS0NnCB1jB4rGkPjmZoQa9wRxjq6UZSgA77lNx2J5zf6t
8b9Pa10MflT9YXvhWF63hWNL5g1TpIUNEBGgKkRkU8N6QQS7R2bXESQD//fxd7ovEKoyqQbgbVah
c2tyU0ZbGE3Wqgr2eWKVA5SivFcOlacj+cxbr47rfebWdIGki+YEBKnOy/iciEGFs+gdT/FNYGUT
RHNJOuhDU9b5+q5wrXEEqb95vRDsMyo76nY1XDBH5cL6G/HFDFq3Svb9nLGJpkDWSPGOIXTnqIkR
90mIPzx5AEuwn17f1OCV4NHcGEOTV+A3BewxxnXPNADDGotpw8Q13y0haoeDj9v1PpgqMkfUdhQB
QjhOkdjhMhhJlvQihrz1BAawx3/jIBYiN1N6DdFlPmtdu2K+UELrGYPrGLifyBd4MzJWpEl9Uy9l
45Q4DRFmSqW7EdZQySxrT2m5CQl0xFufzb3k1gN07EsQ85+T6rIYCFeaiok/fisbUH+QzeS3wL7e
dx0Cut9gfZ6+olCv6qCRQd++y0VxIdzNw4hxZeKM0fe/lKcAMW5wRqmzSvvYwVCibKJ+Exyj7lr/
NPUyh1lOGVGovmhroFsFQRJ7CJT2LhG99ruqIJgG7f/exOoKtaWt/4iauSczydpNuOw2cqJQhG4L
D5azycN62xIToda75Zja7r2FVS1KurmLtfedrh2Iam0XCndL49m1PqtB15QWx0zEjP2n/6DI+Mk+
WKsaTie2zIh6SLM42dEKKsJJ4+B8MK/0rUWJkvgQB04xKMw9TRE9XxDmYH1F1/xJqnVZf8T8dDCa
szMhosHYH1pAuyRYaxLUSbqhWYUuxM/RPikfi5fQP1Za7zyVnZp0+P8Cfz7FymPRsxmHcGKSa7tW
VuRYTdOpI0/tBb0sUMnglKokXDFnWkbA/quHnr7t8yZQUkcpL8uUSFsAtcsoUF2f/QHXMFjST5zb
G+0qrzxXYj3JpCYQuJnEoZkzjdXxuLGpDZVdn3m/Iu36J/DPg8QqP0Eoo4TIAfeB2SeraXHZGVxU
bbyl/Ex197C0PYZQ9lyTNeNmLYyGxraXhhX8UK03dfHF/NOqKJETtrNftNfx8kKi8CMFoCcRXT2N
agqpFVTOhrDnsFYS5uwpBKrCwvyQZr2ecb2SfH/AaE2XtpsayncxW8tPfPBxoDwSHrGZN1eIEoeL
6uBYpemOJjlPyj8cwDmWIa0X/RxV9qwJXdgdIT0N50362fG+PwzvBhiukv8WO7hxBzhtw1XHW5rs
LzaLUN2TG1kYBpgq3caPluyiF9gQoEb8AQUOdBIrqqssXV54LJILyGpomR1r7K5jp8RdLBbfu4kq
XuqeGsT/tJNG7pMYaT9+YdrKWbmIrOz1cRijlEVXGd8ydWVzzyxlWgakgqLw3WMgdpBD9PBkZP94
a8QQ2uSrqjhl5fq/elbaT2BWBgimcnfvEH3T15uWTzowhTSYu7MSPiKsWqzWyO8uAAazj4uUNh6y
pnTVesy+If0+ElopgGpwTMaKVQuBa9caX1pocC+kcFZ1DklQ4lRtKkNocHaqF28zeN7By4e58ooW
6t1F37R82jXLqXT8deyv6262nTkc6fIWjM0YmqqXVyoOTZEE/e2ggbPYC+NJfh3UpGyJIbni2RKf
VE7b9i0IQwjDP31UK05Oxr9b7dvGK2/cVcT+epZ8K96HI91ILBwUu8Iwis0WqYFc4iRL6B43K98h
XBQUihxCpdfVnOVvNoBsMDjHw0rE48Jxf0ZGXU94R0mFU+8W+9S6qIT7hQMSI6URM0bbXf0whHDI
jhIziRKqe7zHMidPgZq/2n3PS0bNh2KU+hocN6WYBldl8T1NNJaMDtNP/a24EPf0W51KCRqLAHha
dgAR7jA80mx7LSVjF405c6jjdXa/Rz7lzNK5aENMe7/NiJDy65zp7JkLSoWjEqcqGzx8jWVKl1FT
ykGaAafX8CTgV1Bd2M5vJ4IuzSqNUuuM1x9H60OyfWW6AncRvjN92PKmeoz3sTNYTeG4mWyphZEr
Fdh9c2ozbzkFBV9CaN+5SRcuQ/vLIk5jXHmNGncvKGbEK4R2CDcdaZWP5snf3oYqzunjKc92EYb1
/y5094ZmMTmN5b5mOM3GYrD9VNGszLgHmFo3AKgaPI7slBvsQWoAy9TnyCoATt4EpnVeNU60bmNj
XVr6njDFPnOiwtVj+Xe/VYB/dea7lKFxqbtZI7fdEQAq8DOhqLBNqalTbWa5XQ4JJUnKMnm5NSEQ
rOfDQfYBaAoBCRD9wcJzLjG2/23NffzSNdkDw6IOMQo5vbEXk3urmF1EYi+U5z+d5DVPkkCABrf1
7F9MGn62FKio9mQ7R9GOPkHKMvD50qaOQvpqSg9pB0rA+Km9AV4qz97UNatBi0WLvKUbqCnyBHYD
lPNsScVzBYjuOAYFXrB3Fh5YCxl2NacUBNn/nZuB4DxUNy9d4BLQsQgOOB7Adttd5Mm3Yp46BIww
qjqJoa7MWaimFdHUXHh9TCz5p23kBa6quvCuwGVzT6P9P0R2WbCAJPDYL47TthmnzpTiZKZU8XqL
LlU3nQGSazSKj0Gf78Eoa5WyMmzzeTvLPoSYmMAH01CzWIxkCXzb8h2lQPl0K2zZT0KCZN6EUpaN
RMHeU18W27nMVH4PnHJ9IruRGA3kekRAlinzA7HC8aZr7P1g5HDYcJs165IkN3p3/WYf1tzvTspa
q0q9RckgsPcrEGnIbIMF2/lRBE9GHVQAV4Mv692oDqhgrEStxw446ZMbf1HlpORNuOmaix1GLM77
SB4eF7YmUlYtQEHWlp+UqbCjSLu2TrPUEVY4PSYuBjppPkd8qT/xndVEUpccmTCBeWtSif9Lwar4
Rn33QYTff5sNRNxM3u++Wsl9mlfar7pcs8E1480p0raPPWrz7/2UJC4IYMka8AtrovXcu6mRSVf2
86P4iK9FVrwai67VUq857U/HMwXSWXxmacxs3iSwfOBAi47A0cojj7RGq1ckp4YKLaTVDSXUeItw
58QL5BzC/++13hjgLGvT4zF06lROcCTVc1iK+xIOBx0DRCR/nqQsdvr4O4jCPdSL6ItHw8x9ra2c
c5dxqceKUBhcELZYmrlv/ykEYEuJ2O7007RBGe3ZhvIrqaQwWpdlbc8l3pUTsjVD7VC/MPL4epJi
z8hKMOd8PGasvgJu24UR5wn411KkTfG7ygMF7bMLnFA5acDq7rAZNrL4+pNqPWX5SiIwVranmtjh
qg7UF6bY2ucF1K+YO2bAhBgIovBdlnncXIbDKMf+2k3kPpT601d8Ih3b1JYa+PsLFTqSQmwfzXxU
UvdIgsDu20oVvAvtxlGJbCqR6q1yBGV9zAFxyT36ZatQqtpsmtoFKxoa0LO1xdRvKW6W6khoOYDb
gN1vbuj9B2s0VyWhmEeaWFDuqgpKHZhcQyOMwNNzaylTtKKHvzs/2yEi5u+DDk0XgwCoq6B6bQHx
d/KP4YZ8wlzQv5pa4dzK7faIh3LhN/r/mzOCtGtaNTGsxnPt4SR/L0ZVRSbsaq9gHfqmYp63D3SU
0LQvOHwZIG9ZQIDdBHfT6ynJ/MOYXG7+6MI0NzxMVvjyGfNsWFLULBCteN/EUhTcaVRElFZfZxHn
BW8vrBgIfvtWX6lFAT86VN1DsLH65DhwdI3rBmaLRSRs2Sno7LdCy6XH3mZfbIpj9AIsiJ5X67za
XujsOxBDH/uaBnmGdkS9LgGH5Mdd5A6Kkhy+p52Ks8eCp+/Jl3pkhLHXEC/bpJ5SPPR2T+4TZoZO
faqW3GrNWt5qLdKXIi1fAY4Ygs/NQ55b4l5zu3CIVVoIy72TabZnjnWQV3cJf/Rk8+bG8BwmxBk4
YP9k2ORpGXx3tXL7Ya5fOUFjAvu7UQ94pJdj+L15Gk+y4xlj5HBUbLCHy6enw8UCjlhcEEJx5SyQ
CMY7yVTTZKeiZxIisGk1y0VMrGWxfgivOtrf2g+7QmmROpMryIMGLfuS36eSfW8DNBHmEX2BQvYO
F5h/sCsssFSnvjx+A1uwyZe3rpnk4kufxibC9ypy6mPRQqPVuRx5zhcJLYBTo5eidl+U2uc8y60S
nWw7dmwVKuywkkyJzItlO+dLl1O8t99bxzBtQyqDPRrKEz6H/8QhfTdb+73ou9w4HNbh+VDq8kdI
1WSRoVMGXrYWGx0HxtqBBrz/ijrpsbMq7kAehKNVyvRSd666/HwWmta2DgPab6y1FRwvo1TES8s5
0guRI7bU3HuURklr80GsiOoHt8k8BW3X4tfubKqGKzhfCkMAfg57JsmlKR0Q/LOSly/gGY+No/0d
eOCQmCjVnqqnPV/fCH6GEiA87HMmAHUz1T5sF4yvui+RpfHv9aVDroJ/NFb2UTi/b2EGqmCM7Jwj
1mOs/MwldBQBMn/2nfwBjmudwl/RJrS49aeEPfZgwzvJm6Z60eD7AU8LUDVp8K5dieBwtzR6LTK1
UDVaUlhNQCJPg3f/faZ7fvT2A5qieGHzs1l61U8TzZi892U7KMV4vX7Ov1ykAU7g06eLxLwja/b6
t/p0IX14+hLPpaUjFMl1TPd30wBYua4jfdjITGWLHaQbcf18aHGRgCLiBVdR46Wqu1dXAMx7R7lb
ssJ+Mkm6PMTipDwTznwcH30bVNOOzUwvuR1mrnm8zQYZWGOl9x6KgvFSa6kM7e6FfKViyeuPKiM6
aK7mD+WvQllPiBuf0Zkilj3i2vYU4nfCRPOODOtxIVczCcv/vL8sxerXtydOSrOeMlH9ITdKY/bd
RJOT1Et5ABW+SQ93AE3Zg6MxwMj7jejwQ0Bv9fLo1F28BqlBdXPeKnRSFl8KuvVfPQXGtlJ4Vsko
CxewM8UZ4rWCl7mbr5VDO3h3eYUVAzYNZiJ04Q4KtprblcQyMDocht0iEh51umxMP2dNECsgy7Jk
1U/8mu+yoSm4E79YRdVb7JkIyo7sKbwPFgydMV8HZsPiXQcb/qCVO2a0DvIiY7BhFURko1W2HY1t
mm5m1Ajc943VzeRK0Tj7jxq/7TVzymH0e8ZiiT5bk2ez7+IfI9vdVHLL8n0bvWBXoycmh35bWA1v
N9K+Il5Q1vCiYtTn8b01j4PLnwS2juDIdzRCVVcwP4dueQP7aDGTxU8ab11CEQDmxYcKKh2Aa/ml
efieH9x7lYb4YqHYIGYBmDovIzTp1QSroYsv7Kn2I54wLoP5g2Mb7kQiAYR459UeSNcP74hblnfG
/BM9IWIDs67R5EkKDX/D4YlNs6jt27FnpYJPj/3mpeP7kJi4RIKzW1Zx0ZVGilUf6CfsbEThOxYN
4Hjp4tTUxAo6Qq0eRyqiEe+ym2E8SQ187qirXu/ShsUw1wzXL2RFo1cz6OohmETzWA089wJkTId7
DSVM7VY3YK6yOLZWPcrAxlocIIlUWdHbutc8vmMUkvofWcK3ThGWT+IFY7naSSxbPfEHlPghqH1c
ALk5yVRSFrZhGJpG6CwyswQgzl+zqs332qRbDdD8hLoY2ER6314QGCspkISvrn5SEyxCVS1r6Cmc
BezuMTXI1ApErtmm0KOgrDrC4S9EyUbXq4ETz3Mo1xmOT0wlLP3gKoH6tF/kVfPAu5gbv3ZODDp5
dHExmTkHDR7yDk7kxYRNMqv4TXS9XvkXGI3hus0740Qz/mkJqtwAtov1DWZRr2I+BQ7CUQtu8/On
dM7hXjoze+2hErKoL5NG0ugF0VDb19Mqo6PpwmcAtKlBMa60KPTCNgSOjeOTYUr+aEP7x1Xun3Mi
512b1FdBohxEnVQM49w8JDR4BkwAvkFI7u4qCl8owSwV4XHj/csf28eiGoMe6FOQ+wl7bVCanrDX
B1/G75/S1RG0e8NG1xFHESDtXBwn649Rrre/gSScXccb4AjaviFiEF/8YzPte8lFtq78moHgy0E+
0/J8ckNwSXTdCsOlucPlqwTwKHnTZND47xgr4D88Cy6hKprxf5V6EOVC/QpZJjbijXb7zaosCVJ7
Z64TYlAMrOQiuSHrCkx45SPUOFNU96f8R6a0I9gszt45SMkRAvVqxZ4YpFqDX5zDR0EnBL3tvJza
x/TxGxbWyM/I0cSeJ+uu0Fnz+iEQXWihrCUSlZ/KYxwEM2kKdVSHadB2Lm//5S+aC4LFX1SvXz6J
xxw3mGVd0r6IC3bR/Gs78QcQg/dvKm+LKajKnzUMr/7IJSVreU8+Tz2/UrWSdSn6gnJHmkFTWf8V
Ei+xook0f6eBmg8SRSxoDifSztFbtDbSWZr0vMk63EHF4BEBJJbEwdECNC/3br5bh9LDAj+h+w3O
mW5qVYM3OPrY/DCkUuYdk2uBj/h5Oy/npD5hmZP077XzaTlxPyvuBqXrW/PUUFdLPo3GoPmWaxvT
7CsnHyMCWsTbKEeV9SY09JoA4U1A1K9s5sdVaJOI/+GsPmnBeh1G9s3oNR1f3xQM1KrfjLTHtuOc
B1IiqYaqVkqBaAWPHRBh1Ye5FcwuhrBwu4KpMMG52CWLPbFFJGhFsabFbbsL+AUrKgcatNPHKzhf
VGzU0lqrJUBDKzEPVGt4IIflzd11Z0FS6v7vZlmZ/kxV2JS2UYbvawuZhp1l95pCZtJDtgBA54yk
xAYlca3MzX4DapN2I51MPRClRnxahgoHKMzw6Kb0bszmDGmsgtE50VkWWhegrnvzmB5kQqHe5qPz
t0qgM51IkI0DWLP39yJVYJYphJRGlJqx7CZy+V5Aro/ZZUos/lvN5/+v7HUNIVsqGF+iQKcaXdyc
ipPw1YwZPp3ahL4s0bZ8PUUHDKW1CWImbBPBqcqiu9tU5co3JWpHbQjyrk3D60M7bHLjiUbMscyH
cJTDxQ4QJh1qqg9M46ktkE6R5zamDk0sEppVlKVqJmSEi0AxBpPUhUszVJ17ZVDRC6jKWMbCaAy9
elFcVRmRilWVPQXPAS6GL255wFIOnQJOi+NuQ/fGtna06cXS5hLzvyVA+Ah9QW9mxIq0GROC9Dfa
o0mB0x5DcytkdKzYreFoADJLgZbEw3yFWepJ9F0Ih+igcoTYYDGea0YAXFBEThd3T1Np//UL4gpZ
eZ1rKWp/IpBGb6LJeuRVRF2G+EAtpaK3lsVtAYcxzibkB0t7Iuhv57bQY9o3yuzAGkh914YNNIKC
NaDXL09v5K9+yDbFdI5CJ/1wbHOUTsDxFSFLJsZLwgtvO9EHNZJtAYPzoIa9dcmIULV+B8o0gsDr
IbBZj7ViDB86ezZysBswXqsCscwbid4HfzvsC1JUpbyGzUof2x8G1j5OdhV/bUHqc+8iyhgT82f+
kvcEHZ9BR9s3w+H1MZJSVupqhPGGMW4Bs1GX12bC61J5EgJTbDy9gH38hJj4X8zX7PbIZBG2izwo
Ulr8pQESAXSsngucnK1vedYiSPiZOG8r4IL7AM7vPtgYXRQRovlzQlnKgTpOLZA0gBq6h/Sl2TwI
kUUpTr7iTLYKdjC4gVjXwWd8JLRfL9uOsiB3GYMBmHECDyM58yS2s2x/6CIDaDyA670xMomKjUop
t99+7kPlVw3Z0Hb4Bhjp2zxyHZwCarSM/Ec/2dMRBo2I2e7E2ZdFqBqnh4A10Ctb+9KH/8h74VRA
tTJJFCJcfevAfYluLOh7Ch9KxWyHlsSfH16z54wh56kbkuIDXNispGACtU50fMYg2NzCuQk0tLgY
vrMnS+njcBOzTO4bQDlaGcoGSrPQv+w/topu9aljjJ7azyu193Qq1p2rxiNwEEXXrzyez0PKspOO
ma3hTaUeXOlotIhW/T7dF2Lseq8SFEXkwy6VUVf1IaetZaD/LRjpVJjeirsgpjE0VrZUzg6Szb5j
I8jiNq6Pi+5+YkWYISBL0S5YnbsMUX1HmtKoQ+yOgR1oRa6msQGOswt5Az/iWHzHOi9i+1URY5Zb
SQWCAElc5P0r7GydGX9FSlvH6BJoG45cOc8b9XGvgjcPS08sk2Mn6g1kKhy+hpAgwoJ/GeyPmQF3
J7ILgLZw4eZ08Nb9bit9gV++4H4mzPqhdjwGUlWc8QdX/Gp2T7KpMBVbJCYiBr8lkSc6mNccId0+
itayBuRVlxbKZI2+ndkvDK1awEjzJtOy/wS11rwWe/SFMheB0epBSbjmqj8Hq6+8r3TKecwhAeOg
lHFC2vzkiMRSGV4aL8VIyqIRKNGzfMYfvK2EnqNT8X5gUWM4dDlD98XeZ6zSfUzvkvDNpXhZFelh
ipDcNMWOuAtC+D1TrchuPN1OBWxgXQrOS9rHXjrCNqS3BVwCnaZhjryCCy+cm+nv7a3aJbnUekEm
QOjp1mbz/J6lpmUof/Lgv70kb86FkzTmPmkltpofKRcd3XCTp1i6Kb1bBxvPYtyxXv2dMQtJmW5X
5XOe03Q7kHaNlt3y3bT8Ub4R4AOzN2RzS3fRzW0gQn4ywK3GML3mg1V09rddCdpxpxBLQwj3Z8Co
yGmXFNNLgPPBWep9qzkI/FHq59KZJUE/mv29NArlTR8Gw8kaqmPJ8bLoGyaUDIH4euOWCgHo8icm
yZUrrCCMeznA7TzSXt0nQyWBWMmDcvzVkatgDkUTFATSbsM+5/uBv2rLgocl5buJ/gRRByg757Wb
VMWSX+Qu7D3OSHtkSKdnJM9A9mt2D2PpMfI3wuLYJY3IPgnUCVozKBmVBNSqB3fPmug+Kzr0Xu+F
UhefdFEEzXlVr8DvgByBpW5osff1G44V/DP9l2FOGJKQJqx4Na+BD7XBiRW0P0hfjwbwYEwNJlt0
K9JHa7uV9MGmLB9aKZdL/Ro5B29oWmNXFFED32FS0/lWwVvRBbLXrPzVTSx1Rns0TAOSGlSfvq2W
/a7WoIyzdYsYWwzwcL0Gxb0MccM+A5h1aw4DtmJ//CeL+C1UOMgd0Yx2v0zLtkKzf/trvRlpCaeY
jDAULdKi8iYvgXH4cbqXdDTpP9Ia9OSfVooUhMaN0Tb/cqcstprTTXk3Iyq4Jr2vWrRshSPtDS1h
vmNv4so6aKpTFzU0K0bZJAPidKNUDFVkdfbMqm3Dz+wKKlGvF5PO8o0cuFMFtxyLnFqvO450JWar
pC0Yo+UFYGaPlWd+wcGE0goOxOKAlZ/cpA8H6KXcnBlqcmp8IU3L9+2cPzPvjgDQfRrqPUDZ69Kn
vCvR+EfCJTcL4hdrTDmRp0hymR8fYJ6iADoo3ab38J2NEx1Wl0K4UfIOdj0bOz8fcLvv/ebNpgXL
PlwdvorZtoDASJy6qQUUuEK215XnW0lNCxAeLbujcFhriRH2JqNuxijGzqyPzLEKMEvoudchYjSl
KMmtn/kFCeLZcHtRMoepgIQAL1bVTVLVqXZ38lu5Zze94ShDrIFBzR/+JszhUc5dpG2/SG3Xctjy
o6v6TotgqoqbNSvXYJ3sadFU4BslKLmourEIG2/NFwBMEBYLTnq4foqd+Qrx+Wg+1FvwNqur0bZr
vPUMbL35Pt/p6NiSUGiNXRvZ8zOFinrsJ4bN+Z7krxRicycWiEhxkjmgwgUwsD5DDtXgwmYNO1XY
0zNwmesywIDZIsf3GOX4F6QGLGUtRc3N0RHUazguLObQDRJKWnDDJFD7uebDnqvNEuyySZEWYvRc
SQHd3c5FVrOp6/HtTcK/ewgBQ0fuJ4ue1CxE63uu76Gm8LLqXjnNBwTyFvEVOFNYWZLBgeBZXuaW
mDVlbzrJiHUliF7XKTZP9snfEwW7cVnL2SjwaRx0ma3LDH8peY38jsPv25o3D/COP1pCH4o/iTMw
epj1N0SWdL1ZB3NA4wV14c7SZF3XvCQ6xIn2iDS+9zD6nvqOH0kul7xahBTiCUKVQK3X9/B5OW2O
O1hDC28bKPJRbo3ewSM+R7XoJU0FCR3TZqcdtW6lGB7kzEsQ7b6TtioR74l9fDP+bnpBekAJgn25
w79gmsFi4mGd7uiSFWkQYJKbI4KWDA9vFqIjirUX4v3WFkBrIu8EpWkfxnD1DBvm3+gksUD7AbGS
FHkCyzouucI7pCfwTiPEb+yoY7jnNnlO2rICIVpRel0e3zemgefIlaUsnw5SKv8xhf+98KEGsfRw
LJJ5hbUY/IDdBBgQEgvtTtu9qxD//I9j0QVairrtLD9kpqHsnxrC8Ka0+wlgV0PH9tlj5ArkpIbI
7ALSr2rBmw4LR75WZSBFSTq8a9qxOQTUL1KqG+ckKdJVvOFbLulvUmTEamchVJM0FubvvLHUxfa4
6J4BSAEmdTsW1ZUe+98dW8UZ1r7d5rdsCAEXoolIm1LaHh3vdHpDuVOn4lIQUY66yCd4tv1wZ+k8
NGfiStA3kV75xcgVoqVF3XAx4/W2J0YJ8ERFbiS7zs7vz0rkhEfVE8NZMZdU271MR/3WwVikUB0q
EYPeON5kyIxVdNJsjX4v5VFZ+Dmnwigxj91indS1WvPxvyxBxVxJxNaU2SvKjR6767yXnEG5fKci
FGdcotDjPI6fdlLbVB0h72aVFPgqHRwkq3huXqBd3x+GgjkmC1n0TxmYvToflxLl7b+MEEbB8yhd
DOukz3G7JzgSmQSx0OUpOah3G39WFI9xHnnT6bjx5GmTFvtTsFuohWs2waWT5gRuuUg6dFHTkbSN
vv1KHKqEWGTXVQ8j1VsjbhvjSsgxjO/+xn2gIFacA3d+KopQWrZVGhtZI+Y2MSE2ZJEmQj6TqiZW
MgHiwgaQbmGUIi3BeJ8xPj9m7h3xJaM8FfG9ruXfUyySla6tSRnAOWa3eKIRXad46ta0LpbDF/3d
Fa7/ifOiTlUPSAb18Tj6snTyc2Ai2WZoc0cazlWev+83GjX7APKT6dcTtgHB9bpYlF6AatIvMKE2
OA6TlzPCrJK2r80ibSP/7L0ZRD6xdLSYgL+3S/kVYAJW8iIBPf71hVFMIBWC99oVTiDZGSig6GhQ
5W/GKM6h3aYFSzJiZwHvO5FHjFI592hmEGizbY9WzXvQiJ5PHhJt/H5evZDNBxBrdUw8Z+xc6vAz
jfF5SBuC5y/42vJwdyfcTutRd6G4pw7vljXhnvebpW02la0Hz/DJnshGH7QZDxXqgHRG8FXDgUpn
K3NHUPloDzDX+cEZymwfe8wNJoOpksxFk3wn8pUU+/nnvTOU6mXX4QJXuVdZjPBtp5FTwjpOfMWU
I+QEJ+FSC48PdXlncuVFbaNVzNXmYGM5YwObzQNAhgetAVwPyUcsoChh9xQ3St5op9D1CIBcUyf6
8fZSr9yNwgkGxrqcekVYOgtpUYtITe9plEYz9hH/oMw7O9tYeT59nTR6D3BjTAgXjp9FRQbq+WaP
N79ZmRH1LSkw1WKIMGnpF36nAlsSDa5yn6cdqHDwaX1rLIYZMpDdrrZ9GkpoQW5VYaLftNomP8mX
3R6ztk/hbBhYyx28tU68S/8R8EMYUZUAEpxLzE8Lzfrke4QpztoGXucDzkvp+mDkbQANya00yZyL
CSXLkoqpalNqixmwbezmP+F4j/pMdibJV1LZKC4SOeU0fjy/Ln5sr8yj9agVH97oVqKb7LsQc4+q
SYnsQ5jajtPxGjM7cFR4V0l+ELIkSyV7XcaisqrwqHlTwcapNAbXGPCIMBiU7P65+BlIX5/FB33s
QfP8CxrV4XTecV8heRahFEbRZ5+ossrtCChWTWLNf/Ft7vlrx5LxvPT4y4E4xHSNKO05yhXgWicf
rgCvRlMEQb7Rhp7+8rd0hD2PuaAOxVgBOilHWZnG1A0EFKGbXY1oQ7VKZkWao52raTjWdfpHGDXR
kv8Pt7eCJuhfGJeT6y1gP+02VC86zT2UjRS1HUsLKRmrrC4A2kIANg/WwzMmlv7u/wC7esadQ+4T
5UUz2lTt/KDofWdv9YgddBNR2M8hTHjxXR1hUC0igUT92Iprnyg6d+Fl6Epm3O8PLSktJDnR+ods
NopVwGrN1dURGmt7uSJbe4NwSCdip73Dtnjd+S+4Q2uSVjiX78pmBoKj4YaSwtIVZBvsexd3T1uW
VDOv4UUSgHpTK/Hicph7yS+c5qeOmEVpgjqFc9HVz2oTohXmuxEKSDqxRiWhC6x5TPB4bjh7QXcU
PRnMZ0vhleq9+G9AKzsvM4M886Exk8148666n+K8JfzFPFe3Pv3qApgzXm1MRwVsIlx/0Q+Lbmqc
AJfcKnU9Um4uopIokMtNLNg9ZYP6souEXJX1oF/xS9+jekQCCfW+q5uRvutCuqXYc/YR76EYK7yx
zpT9aRfIt7v6T/r9cyJTYxeRyfGX5ujkF+/B5M/CtwPLRpVgStav+5AY/oO9L3kShGYtda/XpCK2
M/BNtH/KOBtgeI7xVhDM7ZUgm5LgcbV4AZuA9cFIYpyjYfh77gIthPy6iJcev1Rz+sUUfsaoNItn
64p6trZRfPwQ+hRVWK5K/r+P+nTkI5L3tFSJt8aRAuEXFFnXTQ4TcRYEOv9glpHJLZeNBCsqy3t8
uy5du/u4CirIJxWprPFRlWOIC53GLoesDD+EPVm3P2SkYJR4cchIPpndK+AMHOxJ4vXSwb8IKa/6
XnXETRX3ujoubPn7K+SOCIvNfAZJCwxDPXSBLhbmBO5/PteBTifvU0TX1mn1MReat6FgPs6nXawg
9YQSK0SqqCKRhKbRIiX1MLwSCBYqhhXjoZy53+LLZ+bKyJaeEc4M7ZYvUtMnK5MRTEaiyK8M3Knn
95SH4MqShhjX50U+W0HI4cWGUDYP+megFMHdUTYABzrcDAvktSYxWE3LDsVQyBM6uqknwHTnr+5B
avKUz84jNbcfL1KjBlLLbFGsoQl62KU1Am48WFWymSQpnyI86stpTk/te2Ri++BDgbjAEcWLlpMH
n08tZquDp1FVGTdUB9t4OBviLoWI1k92/0bWXNce+bdF3MY33ma4ANoc9s+XGEequ/3wVX0WIB4P
dIixVqNYC7WPrquc4FAQgSJQ5CzRQ2YTxtwrMULLgA6Ko6O9U4w/BSnQfgLOv7r6jsyGMJ8rAWsL
LNpkGERU91Mm6FlqLSNdPHqGChBcp+AVowbEq21wmYhQmzblmmBWMFp1ottkVKxgzl0/u0vvt4Aa
zKDGWguWyz4iZtSA2oIpqItJSzxHZcqQXf2AfEJhj9KeCcOLnsW3U6RYlLjwDpUPwqRIX7Uzn36n
ZM/ad78dyG7RdsEx8RrJ0bYm1kn38xU+jG4jp/y6H0vDPlLJf80z+q2Ow6Wp4dgUQN/T9UJ00oGC
UTPB57+zzolJHGjDYUV6k9vS23t/eoM+y6Nl0c8QdrwobQlPr4SDBSP2dDq/rz8EkCxR4ka1YX0q
kZGKi/5YKBl1bOdA0Fg9es2vnS1mU6qsXoRPcDrLWcjXpHfB/B6TboJx2hy5efFXs3yj2bNXYtXE
l/ArUxRomxFUKnG6u96JSatts1GDZEMM6aGRBgo5JSji19w8ryB29ZBUY+GG5nO7xH6biE/13GR8
H8ckqLzYU6VjRk7RwKttYvb2NKBTE1ijI82gYx9iRtEeSRwDHu24wTzVn7NDi+7ys9/rv/xFjo8p
a8x0fvQ6MYG5XNuQbbgxy7ZlvcDJRoNzCoaWa6FGRjWPdTbL9ipDw5i8v253Opwfm8bJPlJSy0pV
J8cQPXo8SPfZ3vWYtNDFaUQQVRxOmTTS5rtFx47mTVzP7/LOO7eTnCr/U+uQB5k1ZsMx2h+5w6T3
3/xPWkjyCmDPpIRYkLt6u6FXoZmii636rJ2n+aKk0W8/Wrl3sP46I+w8XPsrmcQHw1eUzOvVJm5p
l7ZiIaTqRYgBFgpAe8QXKEVCKo25xzvMJOu/uChjbiARoyfo6teniycBwEypEjhEsNbyVGj2TRxp
hZXRr5QaR4Vz5gzSuYWdm6X/GC9LN3zlAhw5uDugguY/Qiq8qdp0qDBbdkORl9mXvx6EmRzwD6K5
VjfGe7NvAhM9wa+ZIfST36QZzSeEhW2Syz6U8TGA8YtYG9tL3ylIhDkDmUtQt9noxnC3+MqVmqIq
UACsRijy8h+maIihL/JrLNvUDTwL8rqa1+SQMN7gN1h6/z0bWuuIKbyGjxY/IBlqmprm5v1mELNJ
RnJ5l0AIJDfR+y3p5twU7QcQ3RNgTh/zzSEg0oh+3TlXuS18jeb3FSeZ53xU2XfyTJBtlvqOw2K2
D7sJGh+/TG7nEQzoQggkxloSB+/lS2p1SpfsDQVDZrEny211ceN/PZQDsVewwB0JWeSJ4badYFp8
1QJsuY94j4FZOwIJde4m/efs0fA8xJ7ZqKBU7jt2eSgtf4u/mQtEl5cn0bTLRObqdT+oVMNLr4yS
wjONU9j7chJsoL7Ixa04mHwCymBoeBdvr0HXDXYhSuuHeu2oWtZuNtTq5ZTS+Tyz92+TUUzK+y/C
xTg5zUJ2nGPF5SrleBHfHz0byRwqwDVQ4UMjPj7/JyN9OmPQIvy4XN1IQwB+HT4EKadDZjem3II4
VFhz86wtXLw9R1pyqnQUcqQEkWYfCzibANVwT0q++z2PgsrJNZ38xHPZrqghrCyd4d9Zd1WdWekF
1N7rhiV1vSsjMSxLPbTbPHI30GSasFSJf5MECNttrS1K6Xiyd++igCnhThht2AU/vdvJ6vY/M6mj
2tHLzb96qPBQzVejAjmEWpCgCs6Lm8mNMeIUaKzzjTWEM4V8KNagZSpwOeQj/z5pljSI4hxAto81
22dsT1cuqHTLWQadDrQ7BIBjPyz/Eensdkxdkz1Jz7vFXxX0n/YjSLsldt9Qsapl7D042JKKUahZ
MI0VlPG7p+7ZiHHEvTgTgqCcmTZenbWlC9HikfO/qs4CdIFrHZ87bwPo0wSMOIdulm/TYuSIy2XU
+wOUL6zr3CAgIE/nVwH7krsCCNO2xrz/vQJudf13MXVgEpgzYfqAI9mH7IFzkykvNs+4gHMxadHt
Hs06mAOFb8nhVE8jMa+8Tkel3eOfy2F81RRR5EecxOh3ep/jrtAHg/ansxuUcJocHRyjxXY8kXlW
Dy8PbiXM2PwuWPwBsBHqUdTVBiSGJM3NAKQ+bQ/14giruAVva5Tv51cbNJGEPgLxO6tsFIhh7EVk
fCZU6Au9NsmTZW3kBCI6piq/oK/faWsN+aFD5mB+UYqiTdxbkzE7gpYoKQpYgdMT7dj6E5X1syZ2
zN3yPG+xWKwFFz+u964DDmBdIvn+rdt9lchHSMO50ZgtB4V3K8nc7TSNv84mk5HDwnXvHYL/lcZt
QTgwxlsEqsOjp2S0apGmmBpX4RkKcTYShWIzk1oX4uAEZCOG2RTN/fbLyt2pN936H/hOsJhfHDg7
BJc2AN1LqTuMfp/Ihzq2L1Eb86Yfvd6luVFarml2IYS/PW/LAowpeXgtCMJw+ZDnhwqAgyQ7d+QW
K3EmSRUI4lkD2Gt+XrwGMSxYdfakydvx2nyM+6amBqZsbVyiaSg5Wycf1sbPcXqtVZhr/OzWd4Cf
61xFBakXBo7OFK2MTvcgbHvMeOh2BBOWSD38SoLiFj0zjcHE6QLEdFrf6YKDR9d7H65AcBEGeXsG
1i3N3ixkp1PwaGi5tsxS5KaAul+vUFWYpnT3EUaBlnHesaMGDe9S5wbr53BjdAHYNfKgb7vvkSU4
of+A/AO6afBQJZZqVDGeVouseswb2kuWvFpMv6wHgkiBXYcIJ1fIfWQN9Q/BIKcQRTmXD0Hf5FG1
2qiyO6LpubOHHVlbF91R4FTSlEaXMyI0oTj/XIieJb3eisWnb8dTCodEqe7Y0sUASbF37ryHaiku
JpppT9YHOG6kT/OilobhB1wYa9XbUMfv7BJ+AEZaeCnUljUP5Sgd3xtskvytLm8VjB5RM5BlcvjZ
CDhuZg9McCtWuTlYvFn0F/wTXWgZm+6lV4ifdMrvLgl+wqmPSmfYGUSj/8OpL7zybplrOBfm68gX
Ykpc9R3JV1rz5xn6VYW34R3qrrSUV+BwUxuYt6RGdSjvWIuH4G4zXQufZKFjdn1FI8+tnkdPPmLP
gGz3EbHyEkmKYlXC65Vu9QaNp2iaz8kPKTLbQxzAwdwHKqQmfw2jVeG11Batr+106M7Qt4Y/r611
dR7R9X1TFvwVyaCy+K4Nzuhfz27sveUf6mICBgbIkrVhrBbMeGnV/LN1SC728/ziKcQqbM0EyF2y
PRgv5HsSZp6XbJbY0qKalOXc0/0Bp0W++z1Nchd0RWiJAPNaYbVwE6HyHlhyeuhB2Pr0xoEcegN8
z53ET+2+9kTV7czyZM7OnuDGU+CWnXoU5GJrqGP4hpvLHUHN8BK8G3PTtqYeTKXIca0c8VP2ayw+
l+uMeB4EeKKXsgfYYtXx734mj74o/7JMNMyiVX5bgWssZ9pRH5B3YqfNplaun55CmvO5UWenaIdZ
A8rvIEi28EwrHz9Im75RMJmzjJQwgTheVQulvV9Q3ZM/e2PsQJw2rYsOisvyY0Hhhqkqu4K6WBcF
9VONBhqaO+pdyMFak6375gBnD9tTOzknmSiEczR0DxS2nYsDrc6IdD8QjNqYM52zCbtdpflh5Fwe
I2TsCCd8ZpOkzXYwbVPDl9ydDjCesXJTUtT6yHTrPHI4MH57mvAiuyncj513L4ib3kGShf7U+hQo
LvLjiktOzD9Bxp1YxpxRjMIR4WZHsF3pFVexqVjEZCM8JF94g9T0Y4cxWsbeI1y09QqGGQzihgeq
WFA9v8UMuXkJCmrrjcI34lf3tAiuDZei0mSuOvBCf5+TrUnPmrDAKsSCFKhzHjOzhVNxKfZRH0v+
GNkMp/0mWAMX5QFT+2UNWkRssMmJtXx91dnFhjaj0IyJxqIpfNvWVndiCNpr/P6h1LTqcVXKwQMx
TN4ZN6xYvN1pYRngnMIBeKy/VeLTCZ742T0XkpbDm0t3STY7m26ATdA/kIivka6o8usp9P3SRpDA
GXNIh79DQLODM0fcEZJLPUDLag1ZI7K+83eFAEdgwNyeRfrwFTmf06ewM4NjvV3IX0WkexQH4scK
oQxbUJB6Z6F+EMQCxyw0KEKikAPhHUxe8PbXG9Ah6rxIpbDmFaqB9yJAyMYsseS9YNDkfZLXwj3i
fRPDywnVb5JAP2pzYLOCX8KQ4eTgBH71a8iHZLOANtJTgOAD/eqPHBFXrwVMZ7ZQF9UD1qrnmeXn
GQ3UZy3HWsL32eFGvY/NkC44aqayFkVMI9oeAWg2lLI4u/Qhf1rBHQWo4chu3ktJX+5nbruyYF+N
Cvxq2Q83SBf/2ZpTKBXHmRSfVjFJUmdsny2s+z2IpGn9Nq3wxjaFVverPBravk0SdUe6JmJiR2DW
cJJXIElTWcGfE1BnCA0corJBi3a5nUBCqFz13mSBZfM41xZeqeIF1DvdR63shFZcZBE9+Gu/eZ+T
2zmQaajaBvCEmPRBwVbMpqeDHjBRxa/ZAZ+9fz3X0orCkUxIYDYQHCkXVsjrpL92UMvNQbLutOzd
FFPz53zPqBHKTTb+GdZ9VTQ+3TVtC2UsedkRWoOpVyUWYOBTGxGeRlWS63/f5zK8LtCkpwyvzCum
qm5tDM+AkIM0DAfMXTZhA+8HCYhF1KyLbfUNFSC1P1ew5cKs77gPBv2pMxm7RUqLpcgP4seG9JjN
H2iIMzWJNiE6ztc14Hk36751ZhbOkKkKC0NuV/bYwqYF4CVGb0OSZaQpm8u4g6ZrhR/g4YZyOUXc
NzI6dRaArhkJI/NgWNxEU9llr7vT25PQcMWjHKN2aC8N3A0kjLcGWFIjfTTvpdOHj/c2UPJyXKtv
sGi30eI7IWkV/J2guWjWGLv8JxMsuwrKmO2LC59QKkcqEHTX5Ym2A6YtT2o0W2wUC92/2fn1qnfP
iC0gsWwi882RlkF33lhrOlwYVEVP7yw3L3Kx6Gz7DXLPs86YS75rYAIvs1TKPFiXuFDRIPonatiY
lh0I94P8+qJQDl/JbbN2U9hLSMZ8OaNCU4HBOkEizcNW/irdsTx+q4JiFqhsElldbO2XJLrVZ9V5
9zeNy6LANs8OIDB8iVjgRoMvSM38uX2XgcW1wWH6AzyMbzqgKDE3H/21zoN/zijB+ez2evT/sD2C
hENGpvW0EHd8Fv5kbz9JLEhga0Lvzk/ZMtue5/KeK8V3Ucra3tCj9pjmVUfvkKZv1+D9z3gDJo1h
GCaRiSOAfPV9wnYzcFaEVKNeJku8lLSCpXwwR89r/7pLLF+dYiinDY+OKeHyJ2DUbNMW/DPmA3/0
Alvcsxewp22tZSSTHDkeckc3yh0RL7jC7t8Z+whvWUrHNmDBIg5MWVLoEpQYNNJXSVa0V9X/kEvv
DVssR9ufV+aD5b3NPbjxWxbLZHKr9+r7rpItDvBrGgmKvPlcOT8OjIcgZUQIhaYSc/rD5TXwaEgi
uWIEznv11FkdE68BMKIFYn27GQgAKbCFB3z5PJZTD8CQPAJJp4q34fjjz1QtauyL5v6xA37J+smI
4J4C8+V7PiYPgrfNXsn35IGLwx2v3IrTEVd9Pi9VbmF5m4klPxMP7epbRn0XydPWFfBwU3DToFu3
vdAr7IVFIoeo6realqkKAcVwXOHRFFbUeP0Ch2X2iyMRQNjWcSl9BJ0mG4yYR49ZFhC5RY7unMuQ
YfHQZ5E1kDL8r+uI9/Bou3CG2PXE46gYaBB+67VHIdlu4mFGM1N9LLit3QrQ3Ubl80TeucGGOS6Y
pynMY80BtC2RbOWtlDhJw3gBKxaYAOrBn2H1lB+S7SdYgz9xCmf2+3U3hMpb4HJCBuJ5KcZwJ41G
aaOZTkkWOgqTDXciPZ46UGApvVcI6KjW2W3BlQ/9NhLKa3PUL3Q9Gmb5i7GJxZnn7QA3MddF69nR
Sa23ITOETJeaQk5NtysUQeHvPsHHt6fxbCvA5/LSSAhjp09FH1fr1F9n+UiIAdjcAGt9KuNXKSV2
irYQcv8bbVmObRpBIsjgxKFFm1fu4PvRs+Ree+BXbzCJzTxbqNM/aAbLHMSezCCuCrhXqOHOzKpw
Ls/i6uoeNfHBR26KkXuUskkaim8F04dUiQlNjAeivldFoGgwpHfdGmNtIXaPytMvRQGr2XRoER59
3pjHdZK52MpJNQSnfwo9LcUZVJgQXTTOJeVa0x1o62goUNSFwG/1PhkSp6tfKDXI4PyCWPYri8Nj
UGbeupyndoosDq9SjRMhZ4SWuzV5nxZR/rhpfeOAeEDURZT8HKzcYJWLXYBSMZNXhK5xzdgLt/7Y
HrmelBJxhmMFEu0Qb+R5L8f2G9m06M99SGeCsiVbdtYgILBD0HaautCzIKW6ksuzjmhm7PMYh/Wb
ay7GTjKH3Ez3QYx3HUKv2+wRA2uK2M2IbDLyXXfIcqHBfHEfzrA9/QDAM+CWvis/cH6j4/0JX52W
zYjNGZBHnx82Le0pd/KQXx4MbalAK6wROJVjEQeF140xBZqn8X7l9ZX9J0Sf+Jw0gRZROhRb7Sxl
vP0UPKUhOU7B7VkKqEsxEaRuOWlvhPiahpDUmD6Ym//0oKpy33DKLZ40Z0g7epO0b+OSsqA/LIHm
AHXOloN/twS/c/SUV9ChJkloUXiixOpuLM6LwFgimiDeT0DbBbMpmjNWXDUkwEkmgX5hhDv0N7he
L9Z7TJYdTQ/S1bXGnRnBm950BfWJa5Q35HvGMhyJpOc1FoufIunk7xcf2aPVL/F84lE0sS6RDvAs
GpH3vq8Iw0F7hNIw8UOZb8N99sOh/m/twL6JtAxDmKtQY8GpasdgIsSfT/z2kyF60YpXUzXGv6yV
dU+VEtnLDmHRVNsekXqZdrLaM8kkY3wlb5m9W56E3FR1uQU3hGv08sEJgJM5FaJxejHcOeMPhFLC
EEyk16r9buyKHeXBuThIHLuoG8c7ZbQmvjqQDeKxMQrC+bO1nQn3FOFQ/9C3B8627P05bPg4PRxX
mWYYh4zuuIRcfAw6LlZCUapPhYq22Ieim5VB3wrMWIVd5/41rn91c9TiAvvgqZdQc8EuJi8lTzQK
19E52kvDlGabJ9pYVPw119AyR00qPu+nzDrvXQeXiI3GPherd71xYQYRkxLFEHCDiJtebXCa9IeE
S7wn6on2GZvO/3g6piIsK81vpK25icVQIYe+JN/jC5woeP3SISZ2PBnY2uxANmcp8BMn8OK4ZOhw
DpDh1BkzxQ/Bw+rYueHLpaih3u+aiSG0gkfQCkqEga/sgtzzBfX+MxXks4i0MjNRKbX7qFdcv6yK
F4cACQ5l7GnWDTIiqxYI2I+jgXiN5yEvjQFxtgXt+nIL5GGGfKu7TddhmYwqlUiTtbULUHPa6rQo
tYFYxunrZNmzgogFO03/cJBcJws8f0qCJvUCkW9Gt7yQpVbqU9QW19t1YwSLp40BdsTbl5rP5Mhc
vdZhVwoAJzD4D2sK6gAkBWwnAOkjAUUJe2eYMdGTcxK5tmNoCjltpZXXc6Rl44FzxdTMPded52m7
GNCQCIPy0eIeXciqANJe7RTmdrn+nyybIHYicmiC1OusNsZUwBRTGs6PNpauTuCNM/zbymJ7YUKf
QvwN6HvFd0VXuUSEYWxf6i7GVVWNLD5XhA4QXcX+wtP9hiPu76o/lQMIiC5x2FDdTWU1zIevof80
yDxt3zS17cpqSGg9VLvJiaVgF4YY1sdYZN1eh8nbwMjj+/1HZiDXkYVl6oJZiSHhDG8YwVHjDoF8
ZxKJ5KtwfdTrmeZrDd1nyEX/CnsqowVBLGmSfXJBfz3pZ7rmUsXc90tEIEuy+ev2t2DHKCrRYBrG
H75NxGzkoeRK+DFeKdpx2wotxQYZJ4rs4550yi6KB9rkEQznNHpZX+IiD7Ug+n8J06WazP5KdILE
A3ipwCDiskHMqGdDJLS0JN1WdmBTP9lPX04sNLNcW8aVmOcV7kO9Duz1oEp275G1qsAftNuigpnz
DO/ikj442T/c6wc6qIgXQ6iX4EAyadTSx+u2Robiba4xhZ6dgCeEB7FWKIzvaaA4skT0j021NdTg
B7efxDVTBcjY+aNVMRMLY5nzoJtjzHLFg8U1qx29O/5wiE02Y1a4on/UlAcZ73lJCBnXTt55uovM
3TjGh7C9ooYzGNQSXqJwTmAQbAUAXJ/Lzaa0mDVltKro2rAzBCziN9VCKJ1LAMsn7851Zj6hGVwI
s+tIbsNd8C8v767gy83ptaMqNi77GRPl0TtZd937Ub5Zuxb9JwGs5HPXVM4AV7nkXYQHp9U0/O1X
6KM72b01fACTF+zumGTFDYALMGmYMQ5URh5sAFO0ZTsDQKsXpytFGRB09leI4f9pLYCHyz5EEq9i
Wel8kJzdFFexUjIgPonUv/36vvfMcBEjlwk4BoXHbQU+VdfG6b8hNakroi7K1hz0y/HBfVeM1uXM
YLkl7V21SPYBGfb9f62Rf3TcZEcMHJRkCksEtpbUBo3YJG4N2bmwKbdIjNYYqAxY9B4w5KzRzcSh
mLuEkkKnaa+Dk24zSJqzmtA7EjRwL+v4wQUw/CjZlLFLUVVZ7WHm6NQJ9NOLMYJkOx1KKw+l3RgJ
psOnqL2Hfogr49vJ4poZgu3i9CNgsYetY5qNCeJdKuiSnuRo961nj7x31hLKPhF+hx0uZK5Yzu4/
FWQwwUTfA7O8fVOu4cdEHG34p1cyS9qWxFWsKdn/UymRiThrqgjA5s6Eyk9fgMfAj8JaWueMannh
ylbqHZ1R/SbEyydT232n/0IXnDEEKIQLS0GGUu+4FCAGSc1TFuivHMUS0AUEXFAUa8fcjPl90SS1
fP85mzOnNjGm5i88ApAtVuOuKjreu4phZD2rk5wketfuUbeerUNTYDxKX9PoG7TaQAVmpVQOP1Oo
BCp7W7YKMnx7pQzMwAKmEfe0nVg5GmzNmbyr34+LEO8cFPcI4jYGKkp59BPhT3YxgiHLp1wX6cSq
i6+1vGgHtlXZootKJnRsAs+oHR31VOWbYO9YgUIhI5pjB/CTHyW+nFIs+Gy9f82/1cRvzcutTHLA
z0yLIhtOP1doFCExffR9YB9eYBKm0UIexaPiMXQND3/7ds6qeZwQCHp0+Pif2KfL2HlHNNn2LVz4
wnCTC082ahCV2WeSmhEcAjYXY+kmEfTBprMk9fAt4F921mhKR0I1sg0AhrETj6rDZBWdcrtppz71
zxsY1AzL3GhEzpvElrL6y9XBId/+JzZbWYuypAxMiw/X6sKk5EJ605LoJ0M/1vV0WWt3eHV7Q9ym
duUdHgxJsKARmFA9CMAn68ACk7ATMdeG5kgsxQNmAywEftp0N8Fwf8WD/Q+PGRRv3LrzrifIdhKV
PeKvxne0lCY1MrSMipPkbA5rZPqtKfl1b21CpyeD3chdPDUgNA1LfIh4Hv+AnZiqBjeW1fNuLlkB
sBnQ+7jKHf68YhxVccAmcR4Z9g4OyETbI7o65sycpZSWxIBzl/xLAET76cEChJm3YJSbl+A/ZlAa
uUdWhomeZJpsD5UEoVlud0pGahhiG053sDUgcH0bEa55ickuVi+1t/493PAJXihjfj55Lj8ld0LR
x7aUI9QaKAj8pPRq8zSG9nnWVu6dae008Y98Hj4QCM81PwY9QVy7TiCj8GmdFjDufPkvMuUtbGwk
CA3J0mr+PXtNgbLMF9rBJ/SorU6kUnKu5/rPvWChdBmgT1V8n0Yjx1TCtqgH02G6+OpFHgrcNYIG
XEWFg+Cy4/JFccM1NkBsGjLaSUol2nnzutSu6ddTVbpxCTrA8RIqZ1/0ayQ0Q/cexHRhtpMAPEdo
5DoSiih/4CCZPhjimVyqbhlnegoKqHkxcm+WceWHhzofsaxVZLt1JMCzPmFoN0UdaFIRZs40vmxi
x7/CA6TxflydO1Jtk35ism+OGcy3eBhV+XmR4PBu7xOyDf4wG5rH/k0EPP1ZrDxZOWmpgTDaygO9
AUuvvzMELC6ASUT+xbumODL2uuygNrDQAfsXnWuYIkchnc7NgPtwbyPOJgRgrpY5pECZgB1rw5Ts
ssKyM4Nj6ymOGR4/FoHLAy+JYKATO5AjBa0ajilwDdH30uxM7yV8VQvOXaXQIT3W5M4X+E2kRBo8
jabs4RNZldHuf5cFbJp31eSCO29yj5v8t5DlKyF3tTl6yq+EXNg+byKz0PTsDyKLCZxKTHfJfiOw
ikRFNd168/oTa+goXHaxihitCrtoyDBf3far4jYF1TKBSTAZDKBNjaNItOz2BO5WYGpaNo19FAnv
MtpoVppCEHLlfLmSbCeHPoYLFZqt2250EAlL8Qi3Q9oALLl9vegh3DNxCLRAlD/57+lMmd24iPJe
2KsS7EFtetsQu230Jf9S7PKCPHdzV89SqAFfZxGyGG/C4dRaSfLSAH0XmW5pPfaJl0dcNofhkFjA
fXHSUalPNTlkd2Flqos2W+En1iall1EdTrNx7rgQBnycboL8HT9pJ659BiHNADHBKlYrU9zusX57
i2d+5amtfFz8a2m/GK5iWT8I4UNjQ2XZEoK2EdodTYwRFpRXEw7wV0m4qqRFoPMXRGMGQLYs4lrC
68PEmtxd0KNy2d8fO6aqZYGKmChwfOne8Se7e4+EtJz85Yl7K5d8HiHVnaHhDvu/crj8GHZYA5md
jIr4Esth/h04DzRl7Mxu2FD2DnGxd20dB57QST8qvNVBp2xqWWfbTIIEcGWWznh3pNgmGWpjb/8L
lXrn+UBtjuaxZFx1vCED23qwnyPcgfgNIyssudOSgxmr36/sYFG8vBVlP8KB+RugnWgYcQMvwUmy
XXW2gjw2py92SBtgpsiNaIr7YC5zdlDCsqzim1TbgUvX0+O6y0GQn5kF6+Qkf3ZEP0GV0El6sEbA
43fg1XUlq3r4h1Y4IwpgitsADV/sT5XTGCP8C/kNfED5jNOgKOaVPF9DwZ33zHnD3cci0/OUKExK
NBhe1SvtHK0uaRReRJJoz50GQ2Ffo3rRMzq1t0FthLLYRkWNUO/wXSL8rzdzClru3hk/gfzOAmHq
UBssRAyDiONcR0mTsfQHtYmmJCS20Q7qfeQlNwwF/mGEkX9aos0HbgoUNwDy0FSa/2fP3F9k5V95
2FGF5HYqLAOMl/pycfs7a1kGxgH8AC4DxcnruDQJCR+wZZuyN/l+qvMjXDIDKPCrUjal6BYwpMl9
8IzAqqN7goMB4FS+G4OHheGeECLihDT0ympTPAEPpRUkULMd/rO4HyUsd+6rKDWlsHYwSJ/F6jUD
uNl1IU0Zjj6iAxNQB5mjsL5EmXkkQ6LlJ0B8kZ6ZZ26+OadnMr7C/a3BzJvFWqOL+k5AzZjXKPpH
S0QxBOTSIFj4PTWzmxplhmpwI986cuEN2+uOG5o3+Dfi50D3cfOxYNELy/KIJUYSzdlNYq77CilP
3Z/CMCkSI5vi4UNNURuwi59uSVUdqusqAQHwZMCGKIhMPIWBW1n6dd74KPYzlCq+vZ4n9wMJffT6
VRbX3hsk0+o8KqBor/s2Bin03VdDDT2Qcb1lxuWJ7B849PzQb94C7a4kMwq8h3Fhlt1bIZPg5LZc
C6DFHGd0g4uJ1Ze63w1VUcM2lqluHYYf7wsu6YM1lR4c4Na3AdhbYBSzqm2bteBMMNuny3trL3vE
phjDdzW+TbqeT0gzTV1VZR86+n+Aovow7GZUzhs8ILya4di7PpFzaDiyPoWemcg+IPxI/shwbgg3
z9mmlBoxPyViuOXIBhCMn7gEjsyR9YE/3XLH5iNWlYWJMB58TBR6GEQovYRctDS8XApqm0PLubLU
YIc1q0ljgfrCOEyCPEx1VPagLW6pwP3fezGYH5d6PYXqkBgT1ZNnhHhch6bDWt7PLX+LxsbqXjVA
AVKzCHcw6JIbakw+OCC/oVVd0nDGzBO8HExJxyxVczclEFCoWbzU5Pm85Yp/X0GaF6Ef0vSkWOn8
/qFlQkmKI9eCRjXUAud1pNxw+sxYZO9Lly7z2EdvQhfA5Hhj513dWfYWq1S4PUEWCLVmDDH1cJob
DbBt1bEtnvdXB1b0rJUwAS1C8s17fa2iTThX71EcuNwlk5wxy6WDm2/jjaQ6FiAsE692xzeKRnEy
fPHK+k9FzhWX8hfUEbh1Jl24jIz+Wy/7rhuW530Ija12IUNzO669SP2i3MdIyYbfnoGP7ljuBjdk
k1g2NyziJFzHbu499/7zZqRhTRYvg7jiynT52gCFrJA2Qfkb6q8B2cewy/GH6kbCzbFYYeDKqDGh
2ZUeA0A8Zn/YdH6NNt7/rSqd9Av2weajAnK3p7mDKCZLMc4IfGRyi/soidPvdJ4MBL9EjyqYyUaL
CplsohaXOVniUdI8g0y+MvxK6nw6oDI1UUWOEKAkHYgUPybydIlsd6kDKXfQ91FPX7K6kmDu6CfZ
MinykR4vY8LKh9AQ9Qnmr8OKJunMiRP0iPXOUt9XSJtvz1MZ4Xvj627McdzYq3OPQXdm54MeX7B3
mzEc+cbjM0B6QEVZwf8v3fbsrLu2b2KxCmgyYQNZnBNcX+4RWwapr17VD5WXZ++Z5lTebZx5DLj6
/bF0y8CvQQORGnjNN90JdDQo7LkjVABT6RFVg1iOjozcELi/nVOl4dKXXARLnv6Wq8A1Z7m0MvjD
dKQ0vY5qvtWYcDXZUdmVwHfNqa3CdoTPBE4MsOJS+uoRbKoK9Ez4C5owntA3c4yWvA7B1bYFGRkY
GcaiqwfyJZRBZBoskhg9xTnLHsKUxhg/YGExysg0HMLdXg/RqY7scnGGVnV1YcYUiQPvUeML0G+Z
kvwBhxUIdn9Blzw8AHoqn60em4b5tOWwCaHOCQcL5t1ZcdQ1JArxN7QHVd3iHWpUiw3THOuUiE4m
ubT485ZdZG9dVb53BXMBVXKwyqlxiAedQ4A4kKvf91HQBUVQ6og0kO4EyvY3kd6OrGWpVifcw2VB
i2RvENRhFDMUFXZxe9O7kyEy2FjQTXhwGttXQeq4uPrwikNc1Bc8pdVcsi+/4Vs9+jdFxvAdnmse
KR/gve8aOTmKX/S4FQ0T+iR47TW4We4FzW0SM0qmytKA628v1UPGFfvrOWMCcpWOswjj3EhSzvBL
UNx4502cjOzFk2cf9mQHnPb3OdcSg81c0e/kLKleODc97Dxi2N32EehcL/vyqoOOf95nxT+gAgpr
clFUmISOEjZWqQ9V/SEw8VJsxVMXyDELuht9p8375ITlIBWJsbp5Ncy8wHCAJ3/FznJq0M2Fyqjp
ajo8UkAP2CDIb359rEOluurm/sXIWPlZ6hJiz+uQ1aURF5Z7zcqkhb9fanR4+U+be79C/aNWQOAA
8S50B8Faa8iXk0JqSkstbBNcy7I6IKAHhv6UV/DTEVmBQJo6l/Ol2gupL7Tt0DFme1iC1gZiGBOM
/MauEM+46QX8exrsEvYK+OszDgZZSMeKO7qs0FUiEL+MyR+DrcKfjzXreixY+EZm1IoJRvkSpQkP
rem92ZerH6CEqe1juUW7WT8nwA+QWz5yEQuB8WC7i4wnj/gbOBEahas7wtop0WK5bViFC6DHA3S9
78A9GjL+Vd2xOGsEhWzEDcI1lMbvOLLVF7Bhhm36dBwZCDRojVm/qjZuShh/Ll7n9rmozGLLSAv7
Unj2l5aTPQIwlAouSAfv7V4z1T866+qyM7zHVgb/J/ajGpQ/ZAHSfUDtDVvYimM1FErqPxVwHvax
SKhs9iY2A8ftlPZF4xnAIO9thAj0nb9Mm3YXorEUixQKBjmBempXWkrp2vSz1skDg2FVr+w3XMPT
dnLOoMPgmeGk4cmfIFz8eaCV2kW0wBhXY9ohdVoK9Z3extDOAuTRbg+VljzaTjQT3eFGR6R8uiDO
hA9Vn44nm2igk+3lrAx15oGqOiIR1JPv7EksnDm7UJ2gXLBinb/wE5B+lgxsSuuNE7zXzR8M99pv
Hd70hjFUgGOKm6mvGNat+pTjOLNUBxbae+I5cXU19CbSrWRa18crYaU5iz0R9vmj9lI93Tbz9G8Y
W/mTC9yhSXXUHNxTNdMYzZINX/wm6ZoEBKYRhyYtpnGl/JCeJ5ZPYkuZi6rXYoPe7PwBRMW3cLgD
Vwtu8EhDYrYoB8KXyAWoLUnyXLYmH9CSF95WLguRDiK+GP3TNSwpBVDh68OzKrO7UF0zoZcqWS1e
F2BVky7hwFMQU2d0ZxbHpzm7+7v0rib5/7p+Apm5EwENBFBsT2uLBulhvtooHZE07tG1jUrokZoe
P3Xb0OLY+Vt4e0q61N6rcDBsgyZGst+hFlMjWnP7fLDCakuK9c4trljxhb/QACj7bsSE+SRtqLNs
tolqzWbKWZ1YxL+DDwaRuJpXHeCpqjR6HsW/+nDrcmi21AiUkDPUuykiK++vdE3cRKMrQpEKOj5n
hc3yrCBnmm+FhhnuxeY8WSZtWVvIJLOQneSEcIEhJeWHiTqiFzr3yIfMu7s0m3zjeKonuPBF1PnQ
OE6qiZR7kZFqaC8jPgB2/uIPIfPNATmWGc7NeMPP5GEKSLVjs27v1AUIzcGPRL2GoXADiGZGp658
oo3Z/LUraEA8gI75wzOqBJwIaUyuEkb3WD4MwTnmpULmif1wXKjOrBlivJs7hgKTd7OhvW1v4hS2
p/Hf8UyquY3dxb6czM0t8Np31SLZiKHhlbhQLhRUXUBz0CSEbf3yYJH83S7uU94guRjWK8GOMHTA
Pc765MGPNjq/mTHU5MFPEjEKOTHvb042EbLa8EkQG1848mt4uI2uMjp7gA23UY/rkowApdkkWr+Y
J0eClNw4jr6e3NhE5n4qCTmbHz07fzYuCMPL6Olelm9ArG6FrE+KetkfHqo2w3zCoAbua+3JGdR3
5wdAz995DFUJQ4g0cA12SafzRByJWz19626Bmi9fc3Db5dqlJbx6RGNQb29ZaxMEK0BpDH4BzDjT
8hnUeFtrgV37zMlFKB9k9wiOQ2E2A5JfQoGyXhWRBnygOOgnMdUlj0K9lp6An3NWI1jcAp5Brni7
YlWgJy/6xBRLosK5HkdfTjaZPY7sT0hgIkc/yrm7YrJnQA+vtzEppo5AhLFafgb+172qQevYUg+s
P5nGZGDiZJQ7sRowP5WvYT1O2us8qvk9SI5IQI3RYam83Vcx+gFzwyjJ4ouvpbbq7+/bRETMnH/J
TPCbPJhnEqRp3oqJeI2kyHbeIZ4CnJRQlg6/U59gSwRQdYV/fLxk/griUFv35rqxmzGtH8dijffc
tbzhDzKRKFFQti7Hgd5XaOfBYM1+YuvxHdLgK0CjVCl28Q4l3e1jT1fufhGZpSSxMihSSVhZaMWg
nvrjxgLXoNjXtMqqyu4BQiJcu+HdU/JdYwuezG3cfJI3kuP2ujGpPEWDbmd/BhACFdeM2EUWEKTt
AvCW568gm9Z7UTZTxDFkz8kkmxReSuymQkdvnkzA766qgGE/J7JAAMJsdh5PlCTFgR1TGuJ3P5Es
dDgIFsJ74i1Yq/1UNCNqhqsrAohHrcXA91HzUttGoXgtI8EtkQpwZjT3AJO43RAhJOH7h+oTIXKH
iNvxVoCuT/O23Gw2I/byD/K1VlN1mQkfDC2Mf57Nul1293pxVrJoZU1/KxCUjY+uJAG3URudF2lz
k9+s6pFoQxpuFlxX/PKtVER6nxOX41YEX8dB8rf2Tlqe9SQBefO2c4bxZJ0FHY8nxnM9YTVxY00+
B/bK9o56Wf45ab5t1X8MDtrOTv6aX2LmwVuszhi7Zm5JAfyFZTskruoVFfhHfUCR5tAiX6a+isLB
9cD/NQSowoLfeF4yJIHxT5kG9BDXLCLXYhf5/bRgPIGmIPbAxJ+145h69M/e+HdeBqy+znSdaQ0k
KjjuFGRrkLWf9DocsjGtbLIncDuGWwoRzNwmRx0P0BPM7qEVOBJDXUCzH07aG6eY+lgYqGheJCm7
8XQIJ9nEZIMuzsUWMzti4OoUUuLJtU7XS4c7H/8Xu7byqTJ4HcLyUEbIj+3KBLwD9VGvmOgiuFKT
9W8tD3GidX8DS6A5BSpFseRrnKN2B5/QJjYoSjO6/fVlfPAEMOvNI3Ee+5B3EJ0zIUtCEfeTNvQw
A8Xqs4cDroa+VeBEj/11JMZgOxMz1cfMhxC+xO4Akr8Q1uk2uSxNgtBBYoxKutdwU2OjuxSk96Bp
vwH1Z1pa3hsiGiOor0YDITanF4T7FNNNidSOMdA47YEPSJ+jCKUj3WrBdGMaOl96r4aTVA99Xp5H
Vkg6uJeuPH8r3QQhnpgtIhXO3m7kBIyFDi8cE8xqjO9hE9OprlFUqZSBeiLxyEWYKML7jgqofdeQ
ALmiASziK09PoLXVktgT1cWSQI6kYL6r3Ol1B/IAchXDEmuhNJdgAIvN1BrfBw+Yfy4oqgGOBkiZ
e8SqIsVlfr34NLnu0xbd57aL103Bu/q7s/rgGe+Qeh+9ekaHqJyg6RYvDqWlLX9SsYT7vcHKWWTR
KlZV0gJo+RhH62E0MHDOk4w7OSfWV1vWjIozbOF7zScuNpcvtJlsxp636ftCmwQX5VEa2c6wyY8u
N5Co4UDb0jN6RSLNGa8EYW7SsAdfriiJKW0px/BRmopfs8uKJKAhsISc2jkL9jUToaDnuLEfzljo
r3WgTvLlEKmJkvrM1ADEnFIL6ahu0JccJPpPSX8i0kBE+LTG0N+zmQTeGPnVoM5TSMhvpVm+WV1l
TBzC/aO8+NwvgmMLUhIvjv3fahgxb0C4UX38uu2rAhwevWQOVnsju3xH5WD7qRDSs+iR2Z81smP9
Mj+yNicyt2EP8v7gsp2i4OCO5FkOVoqeI+RTIcgAgXfH22HoMb+d7BQCIA2x75Q83i9SxpkcONcs
JguogxTgwtWay10q8HQK7Ofyh3aZNlwqbIBul9z85+Qm+gZMyQdexfMz+vUbu0dfxvSyruYMUfvp
STU4AFxlJJY1kXerrIr3fmtayA/l6nCvSxrJcpPvQ8AsjON1XT0YTxyxMtLsqibniZijycWJl0b7
ajEg7Td7z/CbGmLZ4BiKzpIF7dZwUsl6RqcQWZc/Wwd6AgPwvIMdwu4JITvmlo37rylEYIZjcdhZ
7TFzLdI9kfssQDQeHbOUi7jzV27Ylo9JYE4J5gAoMEEnkaZ9DKhy5B/G+fvjO+3YifL3Rw/FC023
L3pT6Y60aUSIjkB/WjNU8Ao2qV2axtKTQJADd1E+Lhv6PFi3ElPHoQhnxzTlf2jP5zef7s+TdztE
JQreYhabUBZUllrug5Y7J79VcfIOK7q5G9YqiguckEi4htbCYOtv2fYiljM66aYio9QO+UZ6XZUa
cKk3vpP+Sa4MZXqT2xd2lIH0aCofV6Km7xwCjoKm3YXHlNUDBdXse55wAKrtSYfE0+IFr6ETa6lr
7tNxV/Xk8e53vI27lzMC8m/2nESUzlSxUdQD1n9SokDMa4B8kTMQEr48RNnRhrn9ior+0w7piW2j
afBxYXRwaGQ2wG7XgH29dEhgnjepFI+VEyCh9ILE/EQCvg/Km4G5rtkh+G9FdJ6wTNGIK+R+UrNj
XRJbhxZO7t5ZNlO/tlWxkyBxeLB/fl0Bllv3DjKRN0bD1xFL53TsaLquQpONOwP8wymPqZiA6T2n
2sop3ylkVgTDeaiJWUCQzJ/oqeZZKoh/4yt35AAP6YJRYx7yU+camp3IFJ5wTIjgpF7IVjjdhxKo
tCQKplHXm9Va8xxYkS7fP1yPnweYEz78duTbi2V/BGsoApzsgoFotTopEftr5iUiUW2+QQKWpjnP
N1fqrjyIu9My4PAEqENpWfh3xKiVs/EMHqitQlwHLpwzg9jEWriuxfwbDJxNN3vkT7Jxhn1r+hW0
YUY7ne/HXYzurZjYO+6Wn/sgqN0DVTzhSEjKt57D+V9peW21u/mxhOZvcdBlqLY2sJE6CXubq6Iq
6XC6hkNBUHr50kAJ0TPdRmkB1s8PtjgGvJKXlYyLZ+PLteBe4me8Hs6HVlqLnnCCm6lU/ZFQzBrF
mbNJZvwLADX439+OhYnhNL5TQu+NFCWI+uRMYsEVOi6EoQUEDU4F7G40towj+uEfwJx7OrLdc4Vx
Kd+Of08+2Nac4jb8x6FbW39GpIr9NaezOiQH6AeLstncSfS1djqHCeIiSxuLsoKRJMY79iFMurCf
UpB7mxLMjtmH6Mod9+Hz3K8/UiZS9nsJ9NpJUA5r57UAxncnjjbezg9aiR5KSWQ051ZFmodwNDJv
Nlz7MZqN05x2zQrupEfG2TOqMLQOIk+uu1Dcxb+zjFlMiRd13/YufeY48zF9jcXAD7N0UNdHvtVU
AUy8Kipz3VMQHwuS0F9Wxce/WL6NX10YyjnKNVsdUTZvM/VbUkx0GT02aYTYfEkTD0YMDOX9DrZH
4oscltKlUM25NmSYt2jLaydURVyS9Vg4KUAacIyMlZ4JJHdslizqyPb5b589MARmsAw1sDWtZ9Tb
YSx75NV36W5YQN/lqNiEK3MfNf1aK+b+gV0Udvd6GcYMFK224dUGATsZSpPDr2TGGkUxGw56xvI6
meMdIb4mQCnUv5Q8jM+hU8Fo1GDRddqo2jLZ+8R3GmkRSJ46uTanrDRpukK3eplv1MtsMr8KD0mq
1kgRP90wbzX17WGFazrGnZ776FIeLvDOu63r98agdew5Sjg7xtzv3fWTsnKoDGF5VoWeljOqwQ5O
dvAA/1ggzzXg7EQHE0bVaweoMphaw8QmkH3eFjRHKerWJ/I2KDb3lFkJUkjv80KohPENQEOppqqn
IsR5ZItvZl61i6+q6QDDwKrg3IAm2y3TtyR+iJaWmIP8vNrt45Y8mnTImOXRs1O7ZfsAJggT4FOI
NfcMAVbDmPPcLf3IptU2yIGcadJrLf4Eisp6z0S0ssfUWn1Uor+WB2RhNNkfvdTbCuHPkxo370aN
wkWdwONAOEt+yvcyrUwaGK3hw/9IaYRhU7XA/frDrlr3AXuhM4k6Ts3YtzzUtC4IyP9sfGiS6Ik1
ikg5OvsWq3iDIgF4OcSK/ALuzXl8sIC2B2BDugueEZvCuULsaaDCImKjo/tMAbdLPcPQ5OYl9ixB
hUZoK+WdJl7QQV51vyZrCS2kf9eh59yGxnfDr8ry8DbXMqdBFv3UV3EoJUxoO3KoctzW0o8TxUi5
PMG0UmmGu3DXUDWNOtPbs7MtH5tszCJhxAVp2aD5FyYarC02CjGSqeEJJ0Hk80FxX1CEe62iIgRt
i2Y3O5YWdVZ+a0jwj0N+szwCjlrkwuppRRgrJJH2U4NPoRu8X6IGpjZXnrPw+WDoPGqcWrUgSDPS
mb9L3MSIP5+vangdn1I1k7Jba/dpoNa695/dWfzipktU1p8GyluWZ2YWs4clgMRTMeTo9a+WX7b/
LnBcoZ4qv8rpQ41hQAeXRHNvwwl1tyrOupz4XCjfq3fFTWlC1YY4HEx8+i+rneeI19bzm3gcTbFf
zmHx1fT/6tfowUn9z7cAYwMZYbotRRPMqJ+17EHRCCeu84MIgkUtvKevEpgIh26qbHYcjQDAyFKa
pdKgigQpyaMklMj4MuccCWraapLEwvEx/XxYmfB440hd+CQk5UAsoQSEbjojenPMjOKShE6TegcW
02e2T7o3rplwzgrvIkX64epZlCC3kOMcEm0YbaNBN/LZ+wf5JxikwiNuD2B4dhK8yrloLXvO+VBE
rrLtxpdqhM/NSLduoMyipeKtx8G6ITaTTmv/pf0Y1QfooxK/GLyduldfDYdC4FXb8/qgMU4+FdR9
ZD4vQcPuOSSx9/aRJ5l7D/CxB16wMC7EcX7Ans0r6rR4wv9nj7SZoCrTewhiYigw7odltOKvgrA2
BhPoxQ94pkyaC7+9W6E95R2/cI6HsJSug0kv03VsX7bCB6QbB5cplbC3vYUxW5eK24GkohgG4SVF
hMkvZbzpEJHgSkGmreghp3kLeUdFp7LdgoDXcB6i8LuGzAsIpGFFg0GftKtOMsSfvmrk523Lw986
xjtWM8UiCof4yR7A+gcQeN8KA+O9o11M6jR0qzuMaHf9G7BHcFIEYhL33iArZ93ed5MNOtgievnL
a6ECg/G8D8n/AWcingjSlivje8f4pCTblczHEHZgp76wX6WFTM/DYrGyr5sjND0Y82SSK0QhuEOE
64WE+cLCR0wSadV1CsljBpKnjdYdsmvNVrNXTidEn5+MP8tWkwnYPLoy9kEVfPY35HTnu+Xz7PeX
AxrlC7vdKh1eJnzWW5h+KbdVZNCGmNKkaWQNIIBfQ4VYokG/JeEdpcik9qfS4PW192bG2GqJ8Ne3
mmhoQ1pYlieHXgjKFgpqrQeBdWKwRbmLkNvursTJwlzQ2jYu0I55QEAeecTp/nyOAtSOYThqSQ7E
XypkV2IWabXWNNLSC8CFGXV1FelLo/dqrzGYmuAe4rWzDoFqLgzE2sJRKR3kmkQ4YQKbZd3GQmeo
DkseuyWVzEaFwjfArrbDKg0jkYpL9Zjs/bT1Q63lzGPx8ONwF109sWpEcWwCJFz9eibKQmdW5A06
K2xxwL2iuBAd2lS4uoCgPmWluWSgjPdv13fmiPU1j16qqbkqiDlJBCUv3rFtFBkGJrUBHU+9SjVS
ICPRuMdy56259+vuR0UQQZ4mQnnn+OIYAk7RAyWTbi2T3FFX6dgzyy9t3tDmeRWJRuUKP4EJ+W+G
/V42CX3qtx8vOOwzntgqa8J1V86Myomcf+KK6k18prK0uXjIV/LEkl87pL9mdpMM+fguFrgt+cNI
6iIUE8Vzv9hKodI3GTp5OrZqlEytXQaMhg/nxcxU1tB09oPjsvQAaNwjd5ywbQVKqBp6eVgg2KVz
wL0qlHHHsxXI3G096K7QRah9jzeM2cTMK8zdWKWV0mYPIoO8FPseQjYBiIV+dQW4enn9r0o6nlZD
qSlMVBwnC8rhyaqaLqrQVyhRYASc8ZTnbEbiFmaDKH5Vsapy3ObIrPf2f7or937Oa+0ZDo6gxbix
+BQogpDuh37/M3ockAmuHgITHdZKZIMDj4hLDg80se9ExNyhTUl7ymsc9L40R/3uUqOkHVP696vg
tkUxDU+V5VKSO1DNVD4VXO78Sqre55FMFt14Pg+asJFcrI2dDHGgeX5hfQYDCE0dZnJtrSba+vwf
Ut0tWxFfJH7L3oMcmni/jBhHqX62wctHEpBpKjlF04YyLACz3LsQASCnTqQTRTY9JkpK2EUv+Cbm
Uvkb6FwrhnXDuLxkbX8qtJMxt71LYWWEMrEjM2yT3oOBUSuoceBseCKNJ5IUgH4aIgu7hedBtLaO
t8D2ZVYl87v33DeyE/9mPzDx9e8Ho3B7fxytJGcy0lOLpwLh/6Hg6zJdM7nda+gN9VlkOaXTCY6k
yECmjiA4NpM5Ggj36U5zXnWNnwYnhvpMLKrp1pE1khNwtdUOd2KAUOpWjTYuU1Q/E4mD55cR/Wij
/kZXXK9DeUc0GVzWIAGEjQQt+AVHoDg2mg8Oe02XgWftKVI+uJIHh1v0t7uPlB+HM2HX6lrm2V5k
VHZkR80TWJAV+4skOu2Qph/ybmj/fHCypWzXqXvqYgKw8HxAD16pFaoHkrX3hA3WvgrLlSpdA/g2
c2UfVoxdklPwwTw0yqdKXuhU60TITowrYWkLR7mMv691dIUK7J1foi3dp/t5jXq2NcGRG1OgJ7/P
EE+E/faAAdjrKzKJnDlqdPZuhTokiC3RqgqMhudtQ1sIwi7gH6nC9bglO+2klMw2WGxRut+JDuQH
UixVaFfDuaTL8IIHqtY1h5Km2ZfgiCHA2DmqwMUyjRk705BwdI1ytsTNLOppHyIN9V7vtUPLU32l
kOPlXeSEid+Mww+rpbMBkojn7mva7cxRWCUC0YvfGvl6CvoDfd2584w8kQJvTNxhB9ad24MGERe5
VH7IkID5QeeNvETwPUcnnQGpBYh+aiB2fLS9xBL6+FflfLHHpS4hYeLtQpoWcVlgChK8gJiYdQca
FyfjJEUwy9LdqK7LaXLsRslMfNGIDsofY8Oqxs4NuPwBTArjmA92QD6OkNFgFdDGUv6Thi7ba/ME
BhFHG5hi7ORlZQZxVXFAmi+tUSGa7DRSsszWXqMf5Y7hlCEeh66FC1UuPaozpvrzV6bq/ujVgj79
ERYdf3FHlqajDc9xdlT6prEv1H9Wigu4ikFrqNWSOz2TvA5kuH+8x+n8PQ8qmHN4RPUj9rmcyH8K
jOPwMRS/Ce3coV09mNgwSYVA+liUA0jV0le41i7xL15s/2tJ5hCnyuHP595cbpDrdlCpMYnPWz9e
/lf33IRtJuCMNHZXqPSLzIRXpyZJk187f9vriBniNk/uh+dBwDmXgfzw+2eMXsXZu8l+XQn37Kw8
wd0ek3NqBBhukr629ubl+uTVilDHblqZDHBfF4+ke6GIJAZr7jORlSLa/gTHE626AGdrdEulcUOA
1IQ1ZMWeaOMeF57j7RjCe44TVL9bFDiBaRr1ugoTMreh/0/pNjHc+fY9eT09ESfNB0BpJSsLc/aC
LG3ZTje/qXkmdhmITSxgOC03xrGZb4qfQMBsTCPh1SCjGiwUzuwHNSlizcpY9WA/UPZ8/NN/YD/V
B3gxk946lrcVq4cHkYW5iRL/O1gqvFGq6bPF7j2wM+q0AadF2UrMHkBL+CF+28vS2GwWxLdDG5wS
PV6A/fghfi9olmAwidJW0oIxQ0BHBjHv85cYtt9ptuo3nxTnecGL14jg4oBY2XPkjxIL+vNIXdOf
LNc1GHndZxxiT5meanZB/uqdZVhp687ie3O7JN2tcQNjzG6PmB/lln8pmz5iL1XXodTOy0OWLWzH
WIpRuCJkt8G6pG+JZuK6d8+mC0uKE5OYlmI/W7k0xgsBuiIAi61Hl6GPG/SmsffWBfCfMOsRR4pk
bBGIjrZbAVr0MBxth4NbLI1Rfc0CKmpN0AX1YMxax3NKegBlnVz+Xg0xH8G2R9pWkfvoM1UQgYN4
HglssNIJiWAgv1Vnm8gn7JHgJrCLEdtI3zphRJGuEcaXmnRGD/BGAlEpJ4WvvZyOG9TgJWCKpA//
w4BZr2r11F/GB8SNDjXA3WSzhG0a5toOGuT0OyUy7ypzkS888T8HvY+D35/bXVqXzPd/iie4hCT4
KEGmyAjJu6RimvN78uP/bPUpI3eP7Csix1ObFVz1+UDisXSHYozYiDRBD5Rpyh0kOC8YOy22sSlH
2qOfyWlTcq9c8eKzWmQQVZsZGI7T01jiR3jiDCmtbUj/FY70tTsTkQA9fF+ItAH+bWbAGC5yyh4S
dGBcF9N/Ekl7BbtcZtbVXH+jYmmOVEq9fRrzmRn54uQ0hZ+KOi7swiZvBdWsjJvkuab1oqsnsbvu
2cFa5AeGDU0dgnipxcd21+ynU1h1DSxye+HSdsKoJ7IVRLh2Nw16StWoDkNmGu8mgifDSb8nGPS3
WTQfwKHIAiIh1Ybz2m/Ip6H6lCyDtus58zimZg2JZ4PGC3IR0tm/QpvISUHz3X0kQmNRk31XYBAJ
aVsVeHYX/631QGVHwovGEnVJY0rqQOyyMN8bckc703AF2UyxvHoJILomyDfaMee9iKRWsVs/qGjc
QypWCcGiKVtOT5zqv/EWajylDNNt4BdQuwTx93DiZLyLCCsOxzb1Mc/jGBMVpUE3AONCmSzk7hGt
wat873Z9RxGHWRyCQa52AT0z3LupVJIEC67tqL2qU681m/MhtvtTmU47/mG3cEYjJAfkicWanFIO
zer2hvWYnYvsAulCpfZb85FyFycU7Q6xApvGoqprcYpTb9aaXyQx+500rvbOQejQIwO3uLGmJEjw
S0sC7u6mAysZeB+T8BSo7hYi7QyVw50EPiXb5vqYp+1o7MeX3E34x+BcPI/ZlgwmtdZRmvG+rhjV
fvlCRTFlqEoTWb4s34JOGl2d0wxVeD8wBIIcF/fyUxx9S7KKsSZ5GsDUn4Ziy18W91nb73P+siBX
BWjcuqZn1yyWZWLJqoP08BhlPwKq9AjbeXM/VkrB6vygMo882w/x3D2GzKULuzgHlgQIyxE3UFFV
rD6TtPAiB+jY1xY2p4BmAcmp48LodFsis+WT3Cf5A7HajDUaKuCPggJW5+n2dMNAPovk+Dt/JiCz
0mF4hQ3j3DVnkWJ8EsFdTf6fEsYnQRhjbpl6IJdkbOhauCN9F4pAwykzIu2Fr0lpBL/SZNW6l7Na
uStes2nJ/tgCwmvvv/PZfWPJ73igf5gwnF7aHdP/c2DFgUZHpoPCiQsrSn2B3hM+LPHGyPygVz5A
qklaxQZa1gVtN+xRSDW+XGICpEWqjJ6F9WKcw6NEPgJR0lV7Mx406LGIQnW0OcgAtzyPg9Cd/kSJ
CU5qHSOcHXxsl7tvd8Jth3PooYJB78VdWbtrXq0YOhL2BLNCD9PEh5Th9GFUWXGBwtVHPe16Y0iQ
3uaOz7xvn8G+lGD+s+9yGXQ3wS2nnR1TPBzjMGZ8yCW1Nyo7CRGXsfuL8K4+QDT1XlwVc90v4d02
2d/Dx0qGNXkon6dvjVZFf8ra+mpsUBtINb+WSxa3DU992VKpdDfWiP75LY74ci4uum1GHF7BUc/W
GPfWIB93UXx7FukbWDbctU7TsGyBWN+ZJ7//bZ7Ys/fV5WUMEYtLVoMWS9FLtFGkTlOSnO5w8Y8j
tjQF2Sz7yRCu6QW3I8HBpnXz7RWBK33eycZ2T7QjIjDL7Cg84Q3JtgyTZckAl42rsJlLvnZpQtGs
2fUGkEnYRJj6MBsP4nGjGEn6FaxObwXFv8shjAa7Ax0Lza+mfphMOLHyUYsS6WvK3fg5+AyJ2LDS
E1GOJOx9XgWQ7PJwK+0ZoXVxL9cyqtPn0FKSewq6iWgb4ExDAy2dwtdJeMNx9qr7/vCIqpivP4ou
eZwyioMcNDl92gv3WzoX3rPfgf4uFqZC6RqM+C0Hi8zUcxgaSQ+j7c88NxVGPjhKlPkdg0OA9bJm
5FBMMVlYAQEv62+kYwcpTZsMkYuwXG0i8dDedPNCPyweXZ2uKw4eD3SnDL/HE+D9jRDTd3mqSYzt
y2f/p9oq35Eu4KMC83KAniTQ6mMq1v63bVDlISlsvru+1ZkLhx+VOI9gdKSPAPvyqEcrh/kXIBg2
lFyWBjcA2n0HZhgGVn8DrKOU3/SEhFh+/KqyizSfqWb12imxszp6EKVZn2Zro31a1/AAQzxw8Kkx
oJZd3NeBKmAUL7uqNAQUj9lHdwC9m+euE58GBXSJcmgqnqCY4PITjgqBs0xtOzFGPDPfaMu9Vzni
HMDrUD1dGH4IU1OtPRiLagJ0tf4bdGAVXK57e1YjK4N2gJV/YUTs0qkFDFmyjHljPIwFJI9+oY4l
K7OrQi27UWuSL8pevIfDTOofI5zDahMSAG8UmeyUVslAJ/TBFl5fscJgG5KWqL3wex+sX9trWjbN
pcu26byOYyzKDZMlLAkz1L/peJF96Luf+4yumhd/w9rDHZQO6coI8z97bDbFI+xVlMt957WTyWVq
VKwsb95I2ieTmdT6pE/14YtlDr2AHJA++Xd+m+OUL7ac/FQqPMraxW25WAOvOny5XcKVbD9qCAw5
BFIWAjamJzefFZN9xahp3lZwFiHMehHmCd415B4A2UMN4P7UsCZouaq61fmH9j3tIzalNZJNMyy9
pbHFoFnBo1YrgyxrO362cicihEjeGaeQoNMl4RcT0PgURj9N3TEcitUbUdesJhKa4FVWePuES3jt
GoVTI4kbGWLHlL6FmB9szJvY4mPA9xgu85q54zO2Mk8Vb7pmpB0prTAa8MjvBOytxaMHl9kcCk1M
yX3cEOaqjN1k2H3Io2f+DZYz5Y4zkePAzQTg5j1+fGap/+RUC4I5M37VBlhUrmWIIEkpGWVe5UPU
Ax3MG8cFYwZvyvi4+gQNVAFgtJruoZ2lhNvjvJS+RtS4FFP7m/CTBBrnMDwKUAAezGqAsw6TukVk
6RhF8/avpdQV62P92n0PTcAateKM1yj6mOMdOSCnjlJPYb4sXV0+6gL8/TnDB5SyvQITaQAeBgRW
Mt4GX46LLBCQazmA5D5BxckvAoi/4G1+g1M7YylvnSP1vln+jplGgjkAoR9mu8OfwOzKtil8o92N
WtFfBSB6ZTbDBkiNrnZcCDE2v+KSKECpVr/N/bSAhz1X+tCzxmPrNxbcW/AJGif/MNo/VwdYDFqE
zV0UOe8DHoaZmwmiavSMLfbEdN874cOrTYkbA289/104rEVMlm/2vHCDaCAC9+R+sKtPwgsduLOH
NuQWR4yf2rSLcFzMWXL7qattz6Y76vI2d5H9To+ovcySZ2FX+q7xtLf067rgGlLSWro3VgREvShR
sTx5aWcbkhvwx+dURsaPtHhulAWmOeE2BBOrZ/e5ZEHbY58gmxA+LnBYtGcEOAZ9kwntGqB7GBC7
CoMUviQr+MEbQCVMdvAAJI+8A6Rl8BN3dWEoBvz9uWtGNxM8dVR8iez4KPPg5z26UuX1R5FmxKuO
9tD+PS89IkwdCkr2V7MK616pnAE9I11u3890EI8mCGtP6UumM9L7MPEk8P6smy94TiGwtEbXhIYU
0/MkttmSQZpL5HDwxdmxTavjrlojgpuk/OuvuhcJlVpT3Xu3QgmuCToi6KoLRMwz6lDareCsmlcE
0hhSvEttGqApsuvBwnVyJ32S50SOIIPeWAfwR52FQMwq+h4QdIMW58/B3FwXciVEabTSTkkERWGY
LJOGpCv96znj05cC/H81JuxadSNuCCFkHE8WwiFFfnJfMYoMS4WJmXQKwfIi6na5kBRgyGD8i5LZ
NhxfwNdpZaBZKhc6BcizCJ+3iX60LRNNOlZfpbovVv6tszllJaBhWm/3JjHMo8tjofXj++aV5QuD
u+8z8WgpgvRh32hdRrIpSeZQYo+PCP9WzNOaNkRB9ewv+GTiYdpbAJfTRa2iA1IBDJIV/0WwCi9g
/Bh4L80MX2B1VZiMxSLIkUIDyW7ciWK8bkkVniiRpYFqvvwLXKo/T9vSzceVfQRHieWFS8XCp5no
ownTNYJ1Cv2KnvB+XZxxGennC58klOOqVmhXIU/yd2DTTunGW7emk5MQ89x6wPDXdtYfM/q8rLL5
NbspiYn1nwGmvZMXfjHDr2OH3g5PnbMZylV+b5EiTYYs57K57pC0ErKrPw/38uzft8RR2D6WCbOt
AVTf1UcJcopKtQpizQahMOV/UUgzA0AgLHdBMezJ+vbUHce+spx7VNQnoYNX3bAdvBnNvOvaFFDX
LLY1bIwJwgKtVOwiVFymCTrRoF2rAjGsOkNlz4L0f2hXAr7UatexZ26paXzvfKD5cd18Bs1o82Zl
GS/dIcSy3SgX20+VZ59IRfeqjxRNXKBtJkKIOlYRedCDT4WzM6f5MCTJd3+yryP2xCDidWikpvUD
XMI8iw0WLVz7uQzgua4ai4kyGp9Ay+1mDUEHHc3PBiCjl4IAFBB8l1nPsF4OFLrtAmZWbkBxwDBN
gB5/6zEc4ugGjGhvj3GiMHCtq7x+mOaDj+luAUxU2jz86njsVbp77VGJ9aft/YVO7IhKk3pInBGT
qGUgXBqvHuyUych1eU7VyCkbPXfg7veQ+gVU7ThIojtXuRfKAb6HIzDboZ41Gsa5Jw92VMoMA+3i
674cWtxzs7lx0A3OUi/pHshgbp+Majr2+yy0QE8LpySfLB2VvVvZia0latuWzBlKFrkESl1IjIfD
uh0CvkUEoU0DLrMgPVwKkVzPsSfTmSt9QNgp/zsyzJje4dNxzanABFJvGo3ginGSMNEeZE6QcIic
xz/DxqXnLUfnDlsLMJ8sb8m/DrqNMV9lNRZqoRruHSvzhhr2+jZp7nZPOwT7MSx7JcQ9RpTohMPd
9wX+56msB5BudNGZcitUIXz/TTWqnpUj/4JK+nxbfOprGP8JjqV47WG85I+MoYT7bhGzPJ6KBZdT
xSq4DzG+ED2w8Qzc3DaCIP5NxEA+5nIyQbDzujnI/iCL0GzGO50pNjX7m4/HBdrBP+yYgLLZ8QV0
MBTdVR3Ktp4OCp4H/UPcal2HimoKVniF4Q1egS8Wkgl/kG+XiRuJxkugGhBXrSeL0iFPUZZpXeP+
mKC06IWMShdK97gAE/KQJxJpH9Dp/Xg25YPFMrZJarE1drXJlboBHolMn1y7MzBd8tkbb5KJOE43
JuClSk5QsAb/tSWF9K/ZrtDHo2sm8eRq/4onzHtCQWfhsHAJrDX4fiwB904OHlQdROkT5RcLILwn
RvriqLLh5sLkHjAh70SdehF2JKRVBHpX6UTChRI+nzVVSTK0IBOwiPYCugpMchIo++y48dRk8N05
nqMNUvZYyA/6yOeXoXEmR+Szhr1pV/5XhZQXAKkw0lmsUoHhUHfFjWS+yGBqc7M8oezBj4YpJhCp
IWr5pY7Jz3ciGpiJPt5teWqiOQyhIARbPiHspQMg8XvJyZaYtRGjpXbWfFihbXrZcHWZ2QIebj/J
JTVKWqQZIrnqlk0xLtJ+GBTbqso1IYraV6Ap/lWddnPnt7EJJ7TuNXw3/1OFY11iOzOcJz7Jz9Le
5hTN5Jw7kB0TdCT9AE/9wFdBT0Sw2D735OxUeXw9kVwDeg6/M8p/ANRvFERbXk1H1rbe+0Gl9mjp
Y3lVDaZFRy3dkjxTU8cG954PJtlInXpIANurY0pJ9hxOAQ4h3LiDxX340OMAeM4m0w51cYWlgceV
u0JqLjllvheKDtJHL51813/eS/BSDxFtcEtL0FTk9n8zSlSyFZhfkHljbpHBwHcjfPFmAL46poBv
bUf/zn13JNtxFyqtBaLC6SzKvOMghsDtsY3IJ/twEZesVW/UlgWy8WVaV+OZt+YxcJ3nHrxIFeWE
rfO0E9JDdoGyyfdKXCsRj9xi5HXJBS1ETE+OgHXXio9BKYDCIsvGr5if08SQvWF2Jv8MDU6mprTH
r0O6NKQHEeMs06WsB4aTXqa4r5IrItp/e9e1VMKmZ1UQ9YxH7+ItK8AoctM1p7gMK84twuKygsx5
pgyJpssgvH+FC7f+oIHsBZ/VfbVerGLvpGUHEvAojcAuelnFTyEsg12jcDg93PkFpzTzC5ixo7ui
7o/AJHlNfX+i+3oYF0FrpOzW34FbrO6x8e5Sizt11RhbfU8FQmXUhhC0qp0entDDjdk0yAt0ifuu
+cHdTAjhPFok2UbGSC+Z4cnqdDvgoJzezxBJz9iUNJAdEV2FK6NoR3nmiXzgs8CoS5cSv55kthZ3
Ww/OUOeKUUj/bHz6Kzc1wmBU+EXOStpJ1EUPzc0330dFJaXn2U7O6frhMYGxiPEN8g4VBq3TpMAt
ry45qyaccoitOaCJB7dMHY4iuQAfiYGL/pCQJW937spKLSQXiDCUcFVLD27/AfhWqjwEY/qrI9KB
evtkLJ3Y6MyG6BeWfD0Kz1USI3GcI2/8uRD9IWRDKpM6/OStwz8t4taVejjwFHex84emxwpeS18c
XTbvhzuDZ0fwY/+3Ds/4ZErQZ6oiKwrDtSFlFEfEw7WRFKK4134JaWaUewKXXosGh5PN0q0VHQOq
Pu2jEswpUKEsQRPSgE1oGcq2H19zCBzbZ4IyL//dedYu2Trd9fBegSJzn7tNdz4cBHMlqG7wQfW7
QCk/LlPNr7VpCzDaMek/fKLmtrkgp42NuNV9eX4gExp0Z3x3xqV3CydGuIAa0AP04GJh4FGoxr11
neI2RocgyqQd30dzvqi4J9q0l3uJ7ipa4cj5RPzGrrP2NMaiTCIvRswF/jG68ij0lYTcbYvcwdda
cJncFrQk39D0XFWtzklytaVCorX7ytCBMEYAfBaR1cXbiRoXYiL5AR9BYAO0giGri+toxEmhaOFZ
fkCKg9pgScAtZr1RC7aAzjaJARmPek+gl3ZxRhEeoPqWnN/MDUWGyvWvDvisvhhXtCpSOBIr4RqI
Q2pvC8eOTSxlegbKeVYkWPvPEHrDgf0Rvpm4aGIKNzC6Et0UwpsAzShhBZ27AnA5PHcEVuHmS5Pf
EWi9h+n82C3/Ltd4V7W8sq46nGuGPfAao824m03mii6gWNRRup1FTnh3c6uXniVWTmNgjrCeDGWc
BFTpYi+gBSkaakinikUOyaHrtmezovs8hyrSPnIdmBUc/IPaOWTrdPuiBeeZGWA1OR4jL+iq087n
jp+zeD/bsXgsbkOiAhmY6Lug3MqAn2BEOjSgMX1hoDOWEdie0xgumy+IPqJQjaGisFhviWWRBh28
6RFWTVu+QSbzPQCVc8TU2gKOXJN+LxWcsdPbjOfY4keqKuKfovHB//ADUOItZM9jY3/rxSit3zGO
PPaoLI4JFvPGnRaeegycsb9cwzsi9DiVcd3XPzz3EbxNMqQRf6HDm502AyxsS212Z9+ZnSA/0d8t
/zoPZboMigfQ89cwUPmymz/RFK8kr1AcObLSSUNIOlIsgqJ+M5YF01c7rYlDoUk7UPv2sepNRmBF
RmZzzLeNwbKhQwJR4qPCtquoec6ktLvJv0+CssT+5PWrTew2+TGTgIUbm10BlWPT/1P/eiBqB6l9
4lIU29GHKn35zjqmcVxhqBhSGP5+PXOxIqR0EXbxdY7CsCEHmPdM2jHXW/Ql4GHdqjZamrBQuWIz
fVhwz2QC0XTvp5HHvPm3sd+FoBGoGDjd9JT/Jpea+0q5rQDaBhVwU8uoSjElZaEDoaWJKCfdEk9q
8u92+mEHMxD00g0FCNAmzKFc2Xhwuo+Vs0GY1czfDAmhNFq9pWsuRBqfOkNnNPSqHF8iX8KPkY0u
JF0SmEf0rZnGRS8lPBbUlkSm28YKTU28gy/bLYteVPa1EA3kS416USkUVaczi8BuW//evHO7cm0s
oSAHaV3/ejCit/zXNk+EzesEdHlDOrWP3fKlSHM5UmVoOnIq7eKagrjlbcICNC16hFBsmS1T/CXd
BMeJbj+shTR2kl4a8A3wvAq5N+MuO8LrJa3Ga+AaTB4eaCoHE1l58IFjExxucSG2plcBGxf5AcF6
+WmCCkEATIyNH2/AkNp1XFe0zoXF+Y/297b3TDPp7Y6yBj5/jrqHqKKm8eFGBelr75tMNp5rAqaD
2mBGhIdphDIkslnsN80YlGURIjpSJQWXQuXTPpHC8gF5vZEUWwuzp8tJ4jyDYTAairEjJIKhBBv8
Ptwspyh3WV+RbY18lG1XaAgv0ynzczo0U5nJVKJ9ZgXTBXEuowPRUfQbTflF83q+iFrxPDR05ySK
yY3WE3dL5ds3V4BgecyVCcuxTAlxS/X0l/ld2PVCKMko+CNsEUweFx2DzoznCZnD8UBUhFecmSSe
Hfr2BW7DJyaw2LLYmKid0r3kyJfmez5qWvmnC2e3eu01BBYHOfjkbUYQSFnzX1G+czUTgW83HFLt
sg/n4JpKS2RXms6Pmtzu559iBm54TfBqOTAonYgRRCA3zZPWzi5kyOa/LSe3vNEBktSkgzGyhP4Y
2jHoKBJEcmeqtAvDdEaeHd97+3K6/RciDCcaw/idSif6cDL+GdQg1yh0zzhvPFVyKEZwS8GZx6Fw
sbleG7VXUbxS9CgPHU2TB1qJBuz3O/zzfjIjqYV/MCeMvAWmEw3G83bH87l/GFxV0Ei0BFcroGAi
3pZRt7dxUDctjKhhR9QJ2oHzRX4+LdhbzvJh3fnAOjfqvGYLTQvUIjDqPc+jRCxdxcbC1+j+hdkz
HtwYKEcPkJoVDI8KqWH1ZYDR9Aj1GyxwkjI9l3EJjAnGXbykM3j2PCVisMomn0tgAxA2Sg93k7GO
xyG/zhY2pQN0Fwm5r0ZkFTJA9tXBsvY1iTngBL84TEBvwqUo7NLjSJgE7Yeyo+vIQGEt82acNZqj
a9fPwbnqLVzbtIKcX9CPhXcp7hOjceT8NDEoCVXCxG7fQ6pOqwENW2vBLJYIRwr+aMMS3kq90xF1
NFeInJFKzeA1sjGIz20iQMr0O+JrsfeWUK5vbDvoFFAIzEgP4kX2UN8Tr5dYXOfp2nmqsBWcsdXN
467YUhBmJ07SqPcCxVKNMRF+bL4WYa0y+qYnCz8gfXmGFgpnpMYBJFMZ0xEz6QMmme2Zr4n4/jzY
3KFoeaW6DZonwQTYgie8K/a8iMencZRhSHcde0eXgMGj2Oe6QYHPClO1vwOhi+wPQAILxlMkZr4D
y7NZd42+e/rghs0bjiwWXWlmHfSrMe/hisrnFXsAhxbhcPlVb6vhJ5j8EG+TYth3wxYSMY/cyQZx
ajgULWNBatbE8LvqsccCapkbZkZBZIwQf09B1BziMUvwODtzRTRKpMX2180nXrIS/bKqmpxIt4ju
Lrv6usdo5QCB7rSQTW+MbYPwSoQ1BM1CePcbPNPMEVngsGbwYjrjGGlLqXx9vJ8lD19rTJbA6V3y
ZOR/5f7+tYR2z93GZFqI3boTeoU+0NzcfEvNbg9jzbMiyowkc5XzalNh4d5Cb+1Un3vHREqPoLyw
vC0cuoZteJ1weF4S/F+4uFDG9OEGcFTo+rvCUncuDjJveksqhUYwI6npP86QbyBiMyVcM0EAyxMM
RWcRGiOWMHrXKhtpWDVnyCNp0kXNcb6wA+Nr7NN6K9IHsDArVQX3IweL4eWA/Vo0vsrH1wxhixWJ
9jhHS3uWAJOP484uoW+Y/i9/3Fhb0S+YeucMCy79Owel2cMwBHOtD8kf7ipqQnLIBMwNB+wN7K4+
DcR5VeDuX7TWrtbBvn6UiOKWvU/uvQpWfjqmsX39dVhcJRa2nGEwPdyS2lcPlmTpp2FGLtXgFaMW
4ombVDTTsGAoHbRaZ3xICAsyqQqvAlxMHEi58/NvtM1G53UoGTkrcIdSgWo/po2RwhTEt3KN+FE6
1J38xpSPJOzjMymcl85+8f8ftsqk83IQHf22Zvnvhx/mceC+3hk6SogAP/U5aZf0mmFFteAGaOx0
LT4Fv/dX4VJp6GPnQ1iKvuqjvvk5Y9i0PuBUCkKEK7thsKU5IRks8qr19f2oCLH0n+08K3gQ3Gdw
vtj7tINK4NIq7A5F/BaDXq9qHqsihVDIVBC0iIBch7bvLVSHgB75Xd+lCkO/VA6rgB2MC2XAb+Fp
7q2IHvtv6yT3WAo5on8pU22YWlJ/gI3EkhVpl8mDp9teaFjOoOWIb3vopcgL5d/PlycH3Xhw/aVr
P9WY8uUqZ4ybeP7xNoVJt3aT7TRtPenA5i788nqZ4aEuR8FQB5kC8goIXrqNaY9PZLwn8cyrYDb4
rkM6l5X3z4jRey5yQ27dVHZuRfc9FKpVyjEIffytrNkGIJQuBAQ5qXyWaCK+y/4BWCDUhjAmA+bm
JEEib0DOB1cfFyoLYQH2CRQENkouhzyikd5YhOgvFw3RYoZcal6QZnCat96GqcUvlfWaPS2ZXDPA
bDEd1E9yRTYehEFrtckZltuy9tw79y8wAaRO62hG8Nnoz/2fPlHo6HbDFOuf17HbqkTBaNttrqVM
irG6E7O6o37iOpQFu1loTXit/Ah63YuGmRI8nEXcUvUhBX0pnDz5eVkuyZFjxcjFmSO6ZK8IwkKQ
rRqSXPbxrnh6brT8YQHN6pX+f7vWGeCR8gYLuVhmBPqPo0sgjmK38vCDJe3ZCgGAwKubpOdiFL7P
rwOmIoY7/+avTSVwgkHx0j9lXrqE6GDLvmHQ5K24xjd3/0gyELy0ozIiQE/OC579/koGTOTnQr5p
HP+hHdLTEEDVWOjSiUl3yqDFXmgIHesZPiFDzMA/HvlvRuJgEXw+nEyAeHoMHL3DawtXcDA2gNrM
TEvmXEkSmcRzPzQPs4l+4TKgh4/P7xJ14A1LAvC3FB4hR2mWNo/Pi2VeuYdiwgcWOHgg4buB0prH
G2X9MVop2Sq1n1uDvpv/TVN0MUTlDeo1xdql5X+cwtGD6XP8vIutv11tTe39TjRgxff/jRTbYGgc
m+fYji+0nHo/LYJNFNt2SHHOOXXAbWSHAArvt13/c8qCXHCCcda6ArbxvrWIaLxSb1PG9IJeqLLW
Glo8VClicMbeBXhSOtMY4TfHHujieFhJ/6m/JjLaZHagoZjOdV0lNhq/54f30wmztsN3o3sVBQkS
pNA/yDWE0C5BV+0n6WaPc6Zsz8B7273eyE/hF/lJjEiE/nJ+QzLgs8cRAD81229xYvs4F/zskg+S
nXK2NMnGE+P5Ny9FvZE8TInXA/gg1muSdj1nfIlBHB4MVtbD8OwaxTkZQoEeXxriNJqOes6mTMle
tSk18EdMkOOCLk3Wgu1AbJvUIizYx7jLtmdiFV5lyyuhLDnqymlLcIfoXrS/0krwZAa8vF4ir+PF
zkrkFqRfsi4WYEr25MtNOq8BR1IJaNmuiZLGec9Ks1hgeoqmDR0NxHamEtotVAcLsNkwc37NnkK1
XlOZiqzIOxx75FxqpK33rf+n5ZLS22PwzOrEb4PJ34Y7Ht3YY7qb/tDMMce6GC45YxSBwIyfrSh7
zUB4LMKly2sndW/ShZ9quCBkF+TelJY/aQlY5rQSLmXBlT82QP/dWa1v/VAqPPbSMo9dn2oB/JQt
Nlq8ZEamH6vFLCrWk0pTqjzLLuSHPj+5lWt5csCv3hYs5VMqCExDslDLSfxMO3Se2U68Wlg3M1nj
vyV7+EmWQX0XqrbMJwQszfDBmBelpPma+8PFXqNTU/g+0pFxLeeWLav48oFRy75SriTi/j/j5bXF
gWr/og05Nl6Rn5opFnIdtw9XadjFVp8QlyQyIwiFyc4AY5zBRYHRBIaF4TCEj73BVx4N1n9QaJA5
QQ0a/Q2gF1/8U8hzZpJHYHtBxm6Q3SrxgExhSkGYEzxvJbiq9KXTXqYsYNmdVwnMu0QH6fmptMgw
Fw7wExfnQl3hVvvlmAzM8oPTr2+/UB07ZWvPNzJT4cstACsKFmc7avLv6SKuuqpgwyAFn3Eh5FjD
9IDAoU3MS/M+APArLSnXpjGjZ497Ip/MVRsvqYWCDaAJxFe4eVFAmJyXT3f3PFq2stAhRtMlP5XB
nQoWaDrS4uoE85UbVU9ktaTAsQ5lfg8zj4JmOya4KBzO8jf1A4MWXuEWdhGiN2t88Ab746Rjal7g
06rMkwkYn8Yxz5X7dCNaD1/x7F6iB3vS5ajam6RIv8EiimbygSNMeWD4odR+09sJnippss/hzLRe
mI9gnijJrcwLyQQ4/B9QJTsjI13r3rLi6TjplogCSdbBNV/ddayvoqU2+pzTcKK/tNkPNe3dbkXr
eDqyifve5q8o38QqQnDtCrXGa+4h4gsTGJBJC1yNzVWH5MY2NNBtS6+CvAQSaKgjYpS9Qya+qo2s
bD2yOXXLHqeys3dC/XTqNgjFhpSOwfkd6jBiIWRNBXHElX11MSHAhkAstd+ckF9cm78ZDLmLzYKo
ItDSX74NOxB6syr40PmxkBEXK5wBfX+Ojmt+vobiKQoHj1JsskrCjiO26me6bXj+gfwdaiZsWXiI
ch0z4RX6ZCQofGpD/br3O4iymSihrU9/nlAvLu5fryN9rkE2u852x98SMihRCleedN9NapINPxUQ
SenfEbe35o9wvwMkuEmLwncxRTvI2MFlDPNVhkpJgKVIL+p0lA1p2D7lO3sXZ9VEWGh0m54ovKQZ
BGPI+tFmt4UmRq57DvTRVnT1JNZNJJprvCnhJm6dOD445nfsjjmC+DegJdnW7yrcqXWhgfsiCAvF
+yWWFcDjZQ8zd2hNcfgqxQ3Dj9gC/2SV2FlTfUFrSfwv63VxRjW8CIpDoA0hMNPbiUCwx8WlVUNS
YIpLIf9P1O4LhajEU6beua55Jl1NXuVC2/TFrwvCRJBEBA4Fh8wkCLfcSZY3PefSSid+QB4R/rCt
Lo78AZtdLikA5YMTaHq7RcVs0922dI/BC+AiIH1RJHT9cvrVvI0lG/TlQsn9B2MrAJ3+HF3EbQ7L
q586KFQh+VLZlgasghgwpMJxWS1fjCW8vjnZuxBaKmRHDMkXaUhaMQTHQQYkC0okSzL9/T29Mtnb
50ZUnxtryBh09f7grMuTjqOiKbSGqaPsSDK3/fc51gL8I2GeyDiPHKv70/zNiVJvnt+/lQZCBNRz
UsNymel08swG8f0Lojpmmo6OZQrAq20ThSJ/4EAFr3ESh31P3uVPPrg0SspXXLHxn4EbKszfWT8T
1ioh28eGYYCPIRKbjw2sSJXj9rSK8qQLibWilgMV0GJLBJAwz2p2o7kObqUCGuY2ClYjsmgGQOVL
moExAPfNCmw/xUrCg/LtTG7LhX3fVAbgjihIv7fFCDCHvzR32azFhtvGVH4mcud3DtmN/LErVAaD
M+PYOi0gg3nwimIz6ELCHtZw2myW4FjR5Qpv2GXVS47Va0iEZ/0oetrGHH5Q9LUfoI4NYzc6XXMF
H6jK/0aC5m2HJJWFk25gdY3q1b4SQSMGbZR/4wuq5L8B6wmmAb+lE57Z5cyi2utnHcj3ntKDQ1wk
TSnSm5cQI5QmY3RkAxlHKaxztTYKMo+Uu0Q3Sow6pogu0EYsf6EcdoySsgEDyyGANHrsPAFa4VtL
zoAGZDM4oHv9FHmxu7rpEG8Ov8/VbxWd28KnjznSy5CRb2zr2ylDmoNy3ZZR7WujrdM2GR3Q4xzE
3fgaPug7K8LqJefOMMDVQesStnm2Syrspe6LkCoOdn0dic/M9KVtomgbKuRkScD752s9966vMEs/
z4gUeFLNf09XggF/u3JP0DOvjD8DFhXiKsCY5ykgBsR92Ox7FEOBgNCQwypp+Zi/ombhb2AHhqQF
CMGhaWF4uDMjHKDqJ7qR0d3+n9KKn+fYeWh1pWzM1GBoYsk1XiMErLeQXl0JrFGLLUlVn1iRQqeI
p+Zv11py7VftZWBDntyG0HCLqGUUGeW349iz98TQ2m/rqjOVoEE4iBU54R6wTXs4n3N4qtqKXNaZ
BBKxWj3ER2lJwMv+VvjCTV/TuQ4bPl/+DwIwyG/YxiD8FXXBmSpLiLG9/jQa+NhySQOq1XrhfVUd
eWAfV8DP1cFSCRFN2veld7JNLAPFQqbj/joXsekCfGHZ1w7gZxKtMViznCZIqpdHz+7jGMofEQSh
r41n+YEq4MHmzIaHwtiyoc2OV0iS17V0hc83YtF3JR86QcC/NfswHf8LP78QzhunN5XznYeLa7Ie
MRxnK4Uxk2GdYu4AAlFnpr9YAbJ4MmF2ixhEdYq5YbTes7+lC0V7+tHVnnmY8t9LGPElgHiNvIPP
go48NBb/CYv3n3zgmwJ4EIcMw9IXEMhhA3x0UzNO3oRmeKWIr96KUHLmx/QK6+h+HRDQwAr0g1Fn
RLn/k4CPJ03+VbF7vQATu9H9en+LjSaoXIEOulk5LIKUUEl3mvTmDrf7jPeVLHfozZcFSkeI4NYS
i3mvXffkEUCln/rQLUVPKnmyshrzd2OPME4vgikXvFlxTft3y+ZDkc865sPp3rHHmpBeO4ZTdZu2
3hhE38mZenTEC9GcwdopxjJCeqLNyefKlKQMmFTTd0xQcr8vfOg0t5AcekAqwGwcS+SYspuqveu1
ArhyrZK6W5wNEl6K0F9B1VAT8i084DNay9KdXVbrKC6u/HBz8iq7ITx7013vlV38IlEkCcBvQ728
rzt3by6IHKMo7EPJlKxS+qvTBDIWc1gWTlJmqkg9b4nJcob8qh7Fqe18sYoHMsYTdpWNi2TvtJ4b
dd1w9WwFDcAI4OSI+FDaTLtlM5lkKnUp6W0DbNqmK3Dxr9eNxTC2DPVUc4sbkoYWuOY/lTX7A4we
p55QWFzVB+vQPbYD8cLgVpz09dkkgMZzMIgzQRy1z8IwTnOMkQv9NL2ULEVKuBsE2HI5thnSX7Iv
Uxq8K8H+y/618CCYJ47PXLDbwsL64X8DZo++X3VMtblcv84+JOSt21jaKKdhDXtnBJNnxISTNdFZ
HNt5w3z4GDgDo25LKKPcSiIVBw0KeJ180G7CEE9MjrorppcBkS1f1oEUTzxFdck3gejl2G1C7tFI
6JrG5xhi9S1zmGmYXUxluBSN2qY78mvylRHblnK/wsRmY+irmw/cC+H+X4CAqIqNqNgkydfc1Y4G
pp7zvBHeM+OSoXL6hA4+6hIVAinPaTA04khZNog5WgpHsbdH+38P5mAD9mJiLVRfibhvvoBeNGah
duToqA7Tc0GdbwisaiyODImAtysZVWswpc7NtPHrRlZCpVAFlcaZAreYwyDSdU/vV17iF2TmNdJg
xWO5mjriUVbdm9Q66leub70mQLxD3bTK8pBo9TI60E7hAAoqiE5YkYehMajaHSlUhhc4CqqJFSXT
ECQCTtDiN6Q3aLB26FGwwl1CCmyMCX9G3mpIYXsSBKk0Sw8dorjub48qZboYgL+T1Ezs6zUZcqnw
OCT5b/GQFeuikGc6aiz67+gSUDi4ySWL1kRWMPPlZivZ08Wek2lyWozPmIb22leoUh45Vpo21nnN
xVnhvje0NFmcCyN3f9SYjaDmzQ+vpHxgE1qCINwvedMMtxwtYFQpRMN9TX3ecZFG8oTF58WEdHKU
4XAWzfoFM5yEeEXIJQhqUUEKzx9NzLmWfStpV/dtE2U4A7c/X0wBipNJ0UDlZ9PEJ01Bb3iDlPzG
HAsl0tv76k0dR2T4W3M+7M/j0D9IoP983JYGQu+cn/L6/VyUxD/pO3K8Imj6depEDNwesCDcRVbZ
Ztq4BQ0f/4bEplWzREB5GC7NLJfuBs66/O0xljgVvIm3DlKJQgAURZorOhgDTX96e20w8i2RwkH1
gAroCEX7xuFQ09f8vcxsrHkrHcAWGVdhWdbOEqeMzMUH7SkA0gGQYxYasYCwCL2bwv76tt45F+l/
TqOiqYX8JzzFSj+JPhQ8G6XX/i4SoLWdnxbONLJ4Usi4noU2DmVxlw4XCFK/fM5URnvLEpixepHZ
O43W1us6gbXKLJZ6aHw09TsykedR+YczICO0VB5BJuyxNPOJqIhsdgbtrIk7smAWjrzU7UPEMz33
wcRwHGnvPv7TVBPWGV5j+q+s0fvL9GzntluHRnflpIG8eSsuaUlVErwi+AvT+TbKTYlEs6el8cUd
V/WRd4JhGHRMwHF1gVICvm8OkxBs7ILpcHI3aKqrrt7pIU/1yb2zUFTPH0iA2WVxFcjLKROJeLU3
g++MpLh5dQZ+FYXpH28fBa/tr8SuzXhf5toZ5M5P69bV1YcqngDJbBJPg5Z7A8/03F5eJB5YGbt4
/kO9481LdpKvF7lbmG5xZGvl5pCqpvhBvS/XMbTIDMNqCKgXONg30+VE5hQf/1YnTqimCxHxWaUV
dMO18SrgwO7Al9Nm9DHvQyhJGwlU0aOvvrPgVvD7RNVV1KatAPB2zTF/rvL/WoUCAhCNOElPVVLn
3kYOI0DNq0pqfbXhSiXRZoOqsV4e/uw6pbLDe1ENH0E+rEU5EhkpQS23mrBOZiZxxr7POFbEPc2j
btxzY2UiAHSBZTGu3b+oGcMAHVfVVlezlfSwvDMBaGvSbnprC1y1op1/fDckxACMOWglmqbxj4pC
0UVUOq2M3KJKSLPRdGBWFTokF58pu3K6XbiQG71zl1ESpUv6gTVe1YxGlUKYKXSdVEBy8Ny0Exr5
/NHG3wn0H/8TYAy6SnBN6PMnQOdtd+3XI7L6Q7eRlj6UC0T+xPoTJNKwdTmZyrpBTcvx7Atcz3w4
pQ/vCcdG7bfG8fhhlAH3NEu05DJoWqpc6viQPb7AdU1wJ06pCYhXGwnHW1o0Xo4XapcUkmrz+LHQ
MucMDnMjGZjTHdGh9OiP+7yLhsi3bNLAXXN+Tupd/r8I2gdjadlByUZTz+dYWit59aFTDmQVEkFf
DG9MEvbUU75CMDoc+SpATK2BN+2dGQ4tb7a5iQovfb2tJP0d2DzXkSB2kJp8uyH0hOMBnmG0W0Ks
HXSvKdleeM23fywYOx3dtZ9kstKA/0ntOKmVrdVaaJpd+OlwC5wEq97kcdpajTxXaIOgQbSVi1lT
h9xB/Yfh/2Hbu0Say6C3AqT+YFbR/Vsc612CPSHbaAjxk3n5iM4M7DZ2Vti+pUUnV+NcrCcpoHN+
EyMLiuu7Ns8utd8H9JTUSKpe2XVW6/25XjLRA7lx6ufa8Emh4mtbQ9J3zpJ/z+GcDv5F5RNke2xi
LOSBFFP3RIx1QtowjvKqmvUTol8iEuwOO3WUNHlUv2zEIEWsPQYCZHBO63D/TIb0X5nnCHGX4y6B
HiHflx7hL04ike8Gfby8MpvjE5TH4oD9FV9qAMUjGLRjjWkcYsLNNVzcBkIHEkm//slN/yueYYZQ
myytNxkcZSG4XXKYnB1at0g8++/9+D0Lq4PoHVnm89YoT22031e17j2HcXWpG8j+inUl3n8GuHWY
CjtnsV+UDYFOqmVKF2QhmUoA75F3vd7rHPyGApi7HCz4isnWmIKaJ2cLWwMwxYowk1dddJd3+AC4
widOwaWByJJVstSFbHlgRSoxPxa9UePL0NZkrqBItrWQkZEI/ulcpmk4Lq8HVFemdVymR2EXZGML
OeeOMf+tJ6BIrQIHz9LCp5jZi0HBHHstfVI2l5rGcjDlyR0zixWMJvqahFpmLaXrk4B6e48qpNAy
Z4Osw58O7K0qUr/I3bDyCYgvwskoXcUeENma7pk3NskUVVqTAtlhxD8xoyPvVm3ppkEwn/Cm8uhq
dVMcAFYd0//omKMctmwawA6+uBJvUGF0kgzPvG5k+wruQhnU12HY7gbE7Ar2wE4ZtEeiFOE+eHkF
7uKM9lXDmgrA09mwuSiLQlRfj5U0keYJQPKSP3KK/V+ssE30RZ+eiNaharyd3gKioI5ftSlARM0n
7lOtdm1qDMd6d2VLlB9+LOSdGzfMYDbGJI6N2lNobL8CmjBm9Cp0qoVl3qgzQgDSpDVirS+nZJrq
CLRQhxURJZhvVuY4+ZIjxel+Gwrko69QKJj+Ia92nJHgbT53jOhPkZeR69sGGKjWPIOTAV0w13ZP
VD/Iwup+jRGauy9Z/kW0DRz+h6SwqLNlzv93fYIgNPjUIBT8NovyDu0GaD16sRW3BB4LG71S+WfY
U2wIy4y9iTWx4Sc88CQL0i1UqTr6l3VUAqZcAqmrRN+vxG+az0XqCacu9IDash1hZAyd8D5SBpRL
xI3Ew78yBNNGcHKbt3E/vU9lkOYMxyxsC9EjeklgitmOZ91yyxH4PWhvbgtM8Db23TlAznvvvUTP
zt3Kuiq9wwQen3lxQy3hrGICoOS6JhKY2KVn/N+ox3d6WpGz70OGGlNZxIA7/JEBHbVaTSM70TN7
eonKvFENqFm7f63ELxIrGdJt1rudFk2V2PNO1qqRZqlW0I37AOExhZV5C7UHD5FAguQVbRpjevah
8Fhn5dQujx/EqLa8qNgiCw3fmmOf/KPwnAhI2PltJYKXGGh+cxL+Cl+iU5FzSHajn+crtcMCNVhc
j0ATzmsMp56LyOe84PFoVDiX9ziEKMVNwL/sp+2GweR4lxffU0EQTFuEDjDVbGnrt5gUvSQkaVdC
01GbN7yPBoTEjZqP0otNqTXvflWPHVNItHjWHbUZcL8aMkQZ87SN81i/sXecnAEafflM0NqLWsFT
Y8ILsguBwcq/s+Z75O4HIYWTQ18nxc5VICcEes51vTsUR8FflYi3YHSk5UjQmbLx6ueGv2rtTPhN
Swdns/JimtREVCOMaUa32dJ0CyIab/XF7LLi7kVurqG3t/v/5JoVgriJvscVDusAHRwKzhz0gIqE
OIlIfv7mF8yOyvsqDJitjD36z0oxcG7jL7YE/2sNpms3UpMHDgIZLD6cleKgjRxf1rBRYsrMd/+h
xOJMyrzHDo272z2Cvu125CyLAJgn0C/S9xHyerDlc18ggX+tGPZ7yeLyj6Mwxaunx/HEYScpzNDM
/L6UFC0eSp0ULSFPQNmafmMLQ8KVyEujW6bB2rU+Svm0veymF/Mt4l+hbSF4gr94DbphFO9O9nay
7iylRZ4JaOB5ufVVvva1pOoKZLwEIVCFzTFqDB2Vwvu+pI/0wPRN/0NiA7ugicPZBH2oApHqPoGW
WoDhxpoQx9CU9DbQCrEJ0hDWHXIUulP9TPnIS0XyRK8pSI1YKWlBSGRI7lUHEoz5OW67GOZ7CUXk
Uetoq2eEx8Z3vAo4gJdN0yYYpHwpKGo0iMPxOD0beTLow6yGdIA2Q6OmBjaYnbhCeQYVsGiXkog1
oiUSnjDv2YttNhcAmM9dSZClunK0RnoYReSUxZRPY1jA0QpKq2auV0/Hp9mz5d4gACeRvK0O4DQk
FVdn/OD/VbCTxVJ60myetshefm2nJSI/+oSxKNxSUWMQHQX+OJJhwp9ZdL6LJ1cEJu5+RQ1a7mIx
Mg6z6ZndoZrwk+OZsnySZHOcQ4J0r/gdAf3eCq/rFf8tq6B3KMc+JctrxYqdFpX/NPeyWt3ZM6El
p0KsoTWmjD9mXjVK3gTTLq+lt/bYyEKEzlBeFQ8J0ZZDOcwloAzPM/mEYD3sgiIEGLOs+6xKonrd
pjfGS4y2dy4aUDgHppaAq+aq0ItU4nNeFTc2vRHMtcRX1M5uk4iybWmceEcxKVrYSFnbFz+VwQTN
SRsAthFLrJ70B3NwvgDNL2ufA16nSV9Q9Rqi/jt0KZBC8NZ90NfK+2gGVneL13F49pS6GXALsdXx
GPMe4h0I80n4sUMaj/T2vBXzPiD3x0xcV7G4wK4wfgeTXUb9l41yowlfNGuies/M8wDVPrwYzRsn
cE9FzoYOK7onhxtZBMoXpVwETeUiDBwyoYaLIhJIgfyDHZQuosi4TxAGOAAgBlcyDBoCh1he/oYd
FndsLLumDKd9ceF/lHm/VwhMqpDcn5L7YznuY7eTanW5ScF/VIsFPlXpVC7nPAcNAAncvde4Pq2z
3dbSxKw08GxV0DAEZYK0y9IVoFOsCj/sAOShRLjdh9Z9LyCZbzzE5dkuP3Le3gwbLsWVSRuzYRiE
SLYTeL5FDIg4TQQOswd4xyH2oWwoXz0UbAlRFk7HzuhzpZ3hEvBjRKdHDd0/fCglL8r+mGTUnZ9V
EeCzN4kevAIWLiB/EtreexJfueuO6DJqUoDcNEJ3WKwEtZ6rxsCUIrdUoBBxq5YRAJLyNdXGjB+6
kyi/OfwMYMXU4xKOXvV9TsTBB2fzXZEhIPIVHv9fK2dxZqiRrh3N9Zvp6WuRZMeEyvCK85ztqQxe
FfbuvqJscQbb2imtaCBD5iwjBPiic1ee6Z2eSeKQA2O5yKj2UR/5BfDGaPXBsEj8iJhH4ZhlTiXN
kGJ9F3IVs+aX/Fhqd5vOz4hSju5tBdhfjwEfhUU3JHeGCVz9kOl8RnCCZT8lGxgYs8b5fv/scfxa
kJRu/kC0NqApYRgQwOMcncRIFOvkBaaSV8Cm6rbT6JZ/gXnkfEYUUPQ/eMG/T1RbYcyWJSea1sDK
Pgd2OtLGq90HzOwQlTi/0SGlHMCh74xINmwE1KM6p66J7+M8jUytdR4ndQfCPIgI0Gt1o2vG6GbS
ELEw5iWuotJYpJqhCRBR6ZFk52N6aXEkeZbEGcPS18mZS0BuH4DRf69pmDt5gd6WKB90JEtb6aY0
kXvunYBryvU21LjP1fhX8DhXRi4XIiIbYlShygpTzNDvRS3T8vxlyg0Hg+kvpcI8TqoIx+rNfj3x
ELVwpksgq+2Qq74Gj79AvBDJexWkR2aN7eYbHtaentMB3kn3lGluztq74DFeG//JfRjEfpK2V9Wj
lZqTPf5OlQwKL0qZ5ZX3GiofOKNJJWYMJHNnGK0vx2NRvOc2oA9b6O3zv7fz+gDRf+BSGd9w9nsJ
kVmYKUzyZI2S63INMQZRpJ4mA4TN9siURyz5ByzEuozIX5tDYQgrlmKHYAWUEbIpo/XUloz5/pxt
FKrq3JyeBKO17XKGxnKTZmEXMPtlEsWDXWxFc+LXGAKd0fjhy+7EL045iw5u8O9Qn9wzba/L+NYx
2KGBKEA0uUTym9Nexm52ZXWEfM8ILNAKnkjn8qVUSpr6zF3Z7Qmp5SoKH4IgY/xkGwN9NvYQs9ly
WgK7DNDV05D2EPaXtI4SfyVbm6VB3igo54yJZUEaL8E37wRiAzOmTrFSgOvXFKhXlLLXag0L5twR
qc7kzFNINfMfzmBs7HocNLbOOAMY3rMTI6LHV4AcDfM/hP4OcspUdknTPd46YI5ePM+ZiYhOrs44
ThWcTG1SNaxggr8UjFNzS7TjcjEeoENbasoqNS37h80ge8jEQqwzlNUbpzD/l3Ajwk+jdClnPrBf
9CkzO5EyZLa+vahp/ONr/s3/Db3nTU0juEev4Rfzmm9QflcmnAQ879grM8u0JX9FFVjJ0KW6Qgm8
LsEJmfsVD8VMohGsLhg9ya9xLMvYfYwqGdymKoEu7v6hrCgjNsGD2TxbTfWWA69ibAsnMoWhsK8U
2OEfdx9HlcCI9TciTeDrLayV5ff2d+8JblH/mxPT0XheMrej+e5IxYOgvRhrApCziF/hb/IxrRnH
WX+8SbJ8ejbgynSH4103XpRc1YMPt33uXacTjKv+rbFDyBITeG02JBHypxSTy4rUOWSFQeTP03FM
aY6PGQ+QD6pH5khkzTWLizAZn9DmhQJlJX7ltWYYyu5wweLfmW3YAdu3P5tx9Usu+vg1APN7gsbp
e58h/cjXLAgSvJ0ASta7/tY/RpdfXqJekvXPQVkFUC/bzvJDESMQ9rHhIYipfVuSRQHz3+63ym2C
xb2HQhHHIWHmc4b5gDQDKVnaaRPzYAJ0KvGFfIfh8cJRnFUkTcfnquqZvxSVYFaoeDSxcOvn5CyX
Bm+qyfEoRTcuVoUatMLjOb1Ip087kSVTvmwtLvo34Xi8vEiNnLqZdIq2HXx+z4v1M4Qra+OzA9tz
1v6NTpz6XmivVxxA+EJ2nu2OZujAAKHCqmG7lUJH/1qoCh2LndS+9LHbwtNG3D8LkSXMr6qyli61
h5msDCjdiziSLyGyaJbL8Xuq6k8l+HfOWSvrdw4kUqky2nCD6YamI3Pzm5Ga7Rvs/MgYzrvVsIHL
xzH380OSboPh0b38G+V8vFRMlO2bdBcBujmwDk4g55Nk3CXiQ2EfHKT6fipiV6QiAj877Aelkzzv
IUrjEoB7GAMaBwJZ1ln52F8nz/BEpGP9GHWGh/kIyXMbEPUYLWNo6gtB4oUJJ9zP/sIgtOP+nN38
GGcFCEcg9C4SDFI2XYIby60L+al6Oh4ts72sNlziFJ+4VNWFGnd6Vj3THJ9NkXmz+Y7HTW3QBjWV
M3baX/7Z6zKvHuaLLLFldyFW23TifnU3fHxvTl3xqaMvXPqlaOWzQ8Gj75wIxl0rYtwU0gwY5HUM
aKFYnmUN+z4KAF36DcwbONsvxucS27B1ILqmbRsasYZX2Ewibj29Qs8q61mMLAROORH7XPzUTsZT
yx8BgFWH/ACD23SZDUfmluVL/Pt3HATQeHAz3ZU8N74fqI5DDe0Bhmr/20f6R8uQfWgaKwDExMvD
X/ZdyLFp5vHTVmHM/l1ilbuntwxXh4K80DL0226Pqy+MejTMXp/+9dQjU8dCrQ0uYR5AYAKw9uEq
zid5lgBSUud2EV7G8FYydSUfeZiXrgG2oi0rv02irAZYxW6PunLNGJ9jzDjetPLSwyn6p47f4cyZ
zTxxwH+fO7/bkaljS6F87zS7CRg52+iJiwCjSSL/0LHsFUOpqmHO73RJbQrwM0GmXDZ27IA0lf4k
ormcCykCiC9nikRCpLarn7zgpgBQTUWweVLG+lsXs9vrrV8NuQnkMBwGgRbSBjhPJIVcK+FZtAfq
TqM6Qx+Wh3NHevMcFweMzOnvQE6mpaMye2bbKq0InCfVqXxVtaTd3ZrEdR7/BS6m+MWQm4e7Dote
r72zwS8kZE3A6OQGC8D9qQy/gvgoW7ugoUOpZj7tydg4oYYqDYRw7Kcl6tWvzQgwYqD++FGyzBvt
8fRx1zOEK1H4piWcIeS+i3Zn/6Cn3QWbB63W8pL1POdDUciUdwpUOeC65bQiotWFpGSZNwYfwuzV
Uua55pIZsBvq6ks6SbW1iTeaEdENcVzX6VCB6oqxOCiCwOESzacm+ZwAbwtZcx0YVgm0coaGFgtv
dl3CYuOzwFnVRqILaQg1MTiA87Kk0K956Re3Gsltl/urU1EKnp3dYOqBzMFE2tI9eQAo2/ZzO3XI
YAdsEHrJVYeiJ/52xBvW8YVDDdBCUbg0G04Vvh2U3xbokmO9ZXM+fuPHuqYDJEWRRFl3KvLUbTqy
tyrVtAcf5jGPUxq1L73j34f+ddNC8TGjSKlBmyLZm7eisAOTxy3lxL/i5VHgk98SkOSy07vIrWfR
ewaAl+BJHwwE0rr9Gh0DyxavjjzJ+7mskpBcaxYYW1X5zWugFYv/D6gsSYCVRPjP8eA/r1/tzRyz
qwGfRSj+xX6AW5xTLPwaUwF8+YKCvoZlQKBMgztqFZwq+Unxz8z1TgyWqMc58DfNOaPKxhTznkd7
aVhBbYUPY4tYQfjfeL4Eh2bCWJRD6sJimcDkiGWdFiocovkxypHMP21GdLs0OTETpV526meheGW7
PbZ8/vl4r71w3V5j0WEJcqj+Ibq+jmS2TvCvIAUdYq0LY/XypOv07NKU3u/Ct8wDbuRtoh6MYPRI
Zt+75BBS+YRfBoxZwN9PoB23fhSF7bptuSv++K/3V0XDuib5EXswM2WQtzpYza7H5cmsIacWAVlA
g6Qr7bv/neoRAeNwch06+zzP8Ls6tgqCmMr+dsE/zrCPaHyRaRdzZ/8NNu8jZcc8dLL2Q29A8zC1
n+VcNB1omKKR6+Gs3HChC6oj9R6l5NtuGvOYiw9MqdcZsBrccrhAWLTs36eNvL8miJ49yTX6EVuA
8aUp3cEQYndDdU7R5kFsYj3dOa4+BlBbRFtZiDITvKyVNkR2/z0qntFQWY+tkctaZY6IA+P/S/ez
6Nh9ofPbrr5NoUuw99HxWWMvypZ1r+F7pm3qV73aWxasKVMTjopPjVfHDxPLQMpRFoe6nKJAiQF0
XJtKgTHDoPbftaF948MAL3HwcO9/i5Kuso6gla8BUFGiC2RtDYODp+evqRZnh7S8XsB8ciWAQrab
ZYSpnp/lAiIPAjNKbi2FpODA9uuSoq+ZD49E1pRjdmusY5rICpDL0h4d9CtTBH3pw+aLKQA8w/Uq
yLfIpjcNMebsLZzl/AwXVxvWLrQXHaZIOo5I5JcKwk5ZYdTpG3IqjXVZIBJrlDJPj16K4mFn6Jds
44YVRJW8N4A1kfgqDVfbFcAT0TlM+d45EfkzFZtdOaCD8Kj/Xma9HxB9u0Lj8eG0fbGjdlLI/+bB
Nl3Jx5gR+p9FpOF/h5tA7nBBrleRDBldIs7n1f7oa61Vjz9hoaF313rEpA6p7N/WJ0k01VzsobdL
F+d01qVmnM9JvXV1aXsWmtwKlJFQOeYIttuwQGRY4sRQGFWMIXvNv7xmOMbnC3kprBGjbcossjie
p63riUzeDQ65cOlM4+zDueq87oyP15AqvHbNiDiOn776Hyh41/5XxZPRzvHiFV17fdUchWVEchfQ
nKeh3S9aYAHlrcOgwpEg4s9BpAb9D3zCZUmjskUqafPn62msvNbIovSI+kXLoPcdvaOwY7D3uLsr
Qk5LQPRj0BzujutN9/irdTVzunNulM3/MqDblqfeQsNokB20R0AVsTtcBwz+q7JKz3l6cSaTZH/Z
Q+HL8sqFb935DJDoFKGghJ4vM8ZLt5SBnIE/pGr9FmS81Q/yLlHsSE+SeZSKf4SSO2LeYqzwnaaM
zG6szfuvNgQna5xTOb0b11ue3W8nwsxjn1lViXxoL7MUlJ+z9iRNS4B8+O4/Cqal+4H3f047ARJ4
NqYPecKP/PTxeNVpFJqMGkOoU2Vffn4c2ukg3Z65ZJ+h4IM2cBtvKanmxt/ajoj5W02PAJ1qWLa5
jwxt9Wvt1dVoF41ME6Yc795qzbCv0JhEFU0NKFJ9BK0efGgrZrOa2/zHsj1y+nHZ0RfAYztP5M9k
xs2h1fpEyci8uflF600VFESFIdXyR+8lNj3JVOMChuy0ZBQTDeP3FrvRPC98/490wALgok0i/H3S
YxCp3WLe3Oypzhb2pyUgvTKlhPF76egOG5+TwSvSSuTMRo738o4D2ViCH4Or+mkvRwx3SMaTUaFW
ktnMfeXr2UQRIleTwYW0JhNDDRnlGTjFMbvzyDME+CIkowqSfL2y0+q9bgbKQDmGE8vahNQTxZp5
eljPakpMEGjPUnZaYE6kw+WPJPqN6//d/z5ROCC6CODZ/2olWim2esKYzKTb73thajZH6rtvdj6X
EjcGZmtsfHypCsPrfWvLlhZiF9SpAohYMF/tn/hVEl7/SaJ1V/Y1YywDXwtw38VbAruHtzmw8cpF
LkPPGGWWVzSjQQ7UDeK0nBWRnH7hdyujVae2O8FbAqXLk/+Vke2dqUDzpEf3p/D+sx2NZVIjFbKN
fYIS2xwgvhMzNLqhkBJO/5IryGH5/kLIvfYd/ZvOK9MabXsXpQZXYXno0aSYc66H0zZD1NBzKL1H
uAImAR9kIoiS0n4rIRLjoPnuXRuUuugKcmzS4ZRbuZUfug/9czojDi3LMxeyirf6+kt1byBVcSJ/
d18iBiCdSU83IOtGw4hX3ZtZ7KBrBg9WNxJCu/1Trx6FcbZv4pxn5GRK70aPTzdai5UXDnCJ117h
wayxl9lbTefBgi1VHPtWx8hCsNwi6V5zCVJRJX2QhAzuLCi6Xo3smJ0L7cgrk3S6IADWpFOCFdMr
o8OvKB4zI0Z3jAjUeKWgACyAhEw64m8tAFqP5lNNDMYtiRFrMc6D7lrrYKdEFWilwb3+FPAQHADI
a9VEhc1gNng+ieU56nI6Rm1NRDM/5xNyYIoVirH0LgdqC9PGD18klTpr7nLgGcW9UxORZFshk8a5
FevWpnulH9R9eXLQQk6b9ep90pBB6mxz7r2UEB2CAKE1BJGwfR411gKjJ1qKIhTEIkKBqv6YJ6XI
7fUj/7jDch5HNYaTfyXvzl+wNb/x3e1iRkQvr90ggHcmyPH4h1Wcraqdkq5SFaW4n3XjVu0d2pJx
FoEmCrYaz07QjZfxhPUm2OBjCuj0cfLVt6/SxwivAcMIxtZaubXfNaWGIFCsREFzW0hw5w3T9Xy4
4Egi6GvkjxQC+zFbWSMtfwIEZuC5764E99ePLzGSlNmAZMAxglCczEenn0Zl+4uAPAU9byNFGWyE
uDk/vS1aMCDWtzxKxH/fN+I0gOeiTXjbOgHVi9VHnhGtGiaaJ7Fn0i3zaFeSqq9S2sO09CQtqsm+
o/Tx8ZPygtA98wva3djr8vYpSMam+Y9gd9GqEDTW+WpJny76JxtB0csNT/HQwmQWLaOORQULbod2
eeHwCTdT2+mbxTV201t8wBnQWyu1VJwIkDfwx1O1ii43WglXF2p+fqRkIZJNL67MSzQoujZc39P0
P8kdjqPFwrXCTv5/kOuDDN681gol1J6Wh6SRkRGyn+UwbTa6EjPyi4M0yLm3ficzRpUDRgRU/5Ef
5IDL+5vR1UG0wJNpbuhKTV617k34+U4bP3AMnmSTPnO6C98RYWPCPOVzOfS7IPq4XQDOQD6cDJ/Z
Wnd5/onVkwHzTdo4BOiEZHwWICoyZv0wXNYsrpgRa05BGoJsocKDswC+6hJxlKlcaz55yIfU89Hu
O8rGBXM5qaWyEVXX0poA/MqIPoMxJ+ajuvdesjE9DSJBLBUWpNvfhlpybDOEBV9TqOuWOorpaqeh
XPs4MLFFyiuU7pnUAzshlK/qXjDLrq6dyJgzkOSiCz39ghyyFsAYm1WvNA+koVzqvTLNHzRJCAMJ
rsEVpK1OXB3GfxNyLKurqDr9vTAKWNmD7OkXb7uXxAMQetDGoy3lMCG0zO1T3QgepjAe9TOMZJYz
GOJzjqQqlI++USYgP3C98vrdq67pPvDCHErVg7CrFLaHnEtWQtPLVQ21vugGwKIm4JsK+B/Em1Fm
5PCv92JAMaazEHhnWO2JfcqLLehySC7b0zDVhcOMJLZMrdhrXRoQ+WiP0FrCaXFsKEQ/n1QRdP5m
cywtE+cAVvBp/WrSUcvRknhraKC3iUvm2q08i72HaHwGUiWJJ4qYIHp1sVoRHK2EyiBEo/osXR2h
7V0dkbwcKvqIXQFnnBlhhOsTzqxcWBssgHq+gElCPrDCR0UUIGR4FHd83QKdBjoldzWifIkICDwc
6ybZlo1k+cMgueqa+Tl/6iJufvl2ZjeP+VBYJQbB9zzx9IKnWhvOou66Oa20pvPZQaZlVvU5ZLJx
KWz2C/nojOOkjTEyJq34okbvme/i8JIqzV33XbazrXAtnBcMMe7K7Vnf7DV4apu3iNsnjZH2Bvva
7OKJE3uK0M4oAOlLRdyFyQVmzgxZCoPJT8WPCrfPPHYWX0BlJq8W353IbmntmJYBFn0at7GtHuOa
W9u4AbF+vA85EHISmUduWWSU41JJBu43uNjKm2AcQCeHc+PeZBSrzfHyYIngzzEHyomvo42c8DOT
zR1g61G3eV31zVTEUe6nSJjA4hvnIcmZbdV046sm5m771rmiL30Jjty/2K+53zW8a+xxaRHGeMwK
7lRYPcSNKXPjmb7xNwVBgEr8MoBDIHa5MQEjAYkq1eBDNFrAm5REGGRMM7dqc0hA7aqvaWPi88jB
6Uv6PIzcXLo6tPHXTuf06HPoRONmnFU7yvMpTIPcOoq3pYQJ6rPO1DPzpXFNYEr+YUFR0CgBMIzW
uCmjevb3nX7PKnGs1pav/w1CKSrQMl9Kv4wFiCl/DbWBqZxze7EhT1C3SfG8flANR/HEv/VEb408
wq7WrMgzh8APZL0cIzPfHOX/Zyc84BgFC8G+a9m9p3CPffyw8oOpafvt2blmPz8G2cUUrdDI3xgj
+7EYw51h3faZM4KUyX4lRFNOqtcCulOXytAoNZi6bcgLIufguQbuQiGy8Szh2thWlNgeQDUMVz0n
juBRZyaKtu8vCAE+6T5AbVscY3Hfvs/bvrHHOKDuvzNMT9cBwW8kHk+unxcig7TZrpc/TutzQCDy
lwOLim6EzJ0ngw6qorVMFg9u3/xKCH0mzc667Ant6cx/Krnc3G4da/FQ4hnbjGfht+3MPBKQq1mg
tNsLg1BBXgPs1QdS53f5taJrGSgDZn//HCbB/AYPWZp9JUKteBKeaB524Wd5WTUbm1y7X4AYLrcu
NhOhoBSKWygqmxuH8Roshw9iSwFabrZ1vH+nBJoirDV8U/ReiuaGU/S1Z+v0rFXWodxdtLoUK+Dd
Jweui5pPbsq+U6DcTzRkYXPyhp/dQy9NQdQXhmfJqrICL48WgAAk/TYlrGwEGvw7hVpvzfJmydkC
KBSbpEbcw+EVRm8WsoKVzymzunpgIySmwEIojdbvex+gBLkwK42rjRM2EFfZwHgZDdR7FtegAhti
/p+rOHSl6Ixq47K0FePb9eATdVugz8x5wi3ecxUx5j74YfSmNGJEXdzQaiMg9dMTqVAR/o869233
OVv3ZK++15K68K4nwapOoDd89QmDO9r6DekIn7hVNbKyuOGg9tpwGWXwyozWzOD335tK695XwyDA
nRjU6HjQMjR5YAWxTTKEZqR4kiUxcWqds7DT6Cwd7bcmhDZJNHo8uSdA+26CsoIzdh3fpkaN5fC8
raA6D+P3gZOQr7mLzY4YtvCDPEV7yqkhafV0EqYPejADXMsbw6jvq/Mpqj9hIbVCZWzXypsvK+PG
qL9/2x/OXk6/4cWLsup0Huxbx611cdM3guzLMtM9uIwCDiJLGx87D/M9devU7M0FIQY5XMdjlJA1
vJoqDWsIn1t8t/Wewj2zdQoXf/iJuBdNS8CjgNdikFCPRfBZGKn5OfYzcrVyOjNix+qrs2KnFPBn
o6rm2/I27dQRlrRLYQxbSMPRrvjOJmHcApqT4vQBqKJsGws3v1FPO0gAvGOZN5cpW9wSas2ltKxM
YK7cQ+QXWrgIRJq4yqgDz2+kFlb/CVn2yJoiNGC9j1UoqUgHSIetpY9SLcmBhGed27rweWwyaFxH
zOoFPd1uhYf6W2qfl/zC9Phai4e3R3JaAHneng4HH1R5RlTAEJPuZHUh/ZwWBJBemvkRRvpZig8R
qEFrBarhQD0ezfQlN1/bdmxOAnysthhNPYCxikpK9+1LSE4Px1oRtJPqf5xjKdMh7tqHjzshoCwT
uTyYIqb85oR8YT6Bl+aNWqbszVl/d5n4hQUBBRz0HE8W9QykgPKsuV459LD2R/yWg88DCDkKdGz3
w4txYSipOCrJ3efqxbt3bEQBPQ1bKyzBaBlqvQ4EU1+R4qRsuv48UN/neD8ZGOu7KmEzgNQfRkjf
AVMz4bYOKoX5K6Lzstiv1AjffNJdonHnBu9vVFloEKTQniT0XbSZMQqymUOezZZWMHR++wv6JNlC
UKKObVGbW+47UoTxy/I0265Tctg935+pcHkPKwktLRC9B9p2lDcn9ZqQ4sl8MrLv2TNh4EgILm5R
w0XwxgEfQq8AR56hu5WgHO0Z2vFAJdZ41UHp9XgL74SL2ulLMZiX5R7UwzHTT/B7QHc5OD/s7Tbk
pffDM14rscknULnD6jG1DgDo/tPFQbItyQb1FUrjcyFn2elBA5uZmE7HyCG7QGmDtKKu/4CZJTUr
Mpr9zehMLtfOG54v+++VxCQH/yLeBkSZq0QvJw38DrdyHmw/sonE4TdzhQ2af+iaRrCf5W5TKNzz
sPwBGx6CjK6wxRu97rsNBRAAzVTHuAXxrle4RoTfUXi+jZva446xDO0QXeB9sngXHyChkregMaMA
fzfSD8RTRAhmAso3z0/fjaG4I2at6bsFTV2GnGYoAfkgJ6VbHakoix9+MBDqvxnJKXRGFghR0mTP
GJrFJWW2lx5rb1iAvcV2213zeiv2vvG58ZXHY/uDhoLfaEX8F3IbrvD3Jh3/G13zrCiob9OjMlzd
sOgpr3OylzPbK4F73qYNfbypiGBjGfwYQrHZNV0WHudx+Fe0yGKUTv7egIoCy600LIxhpjAnYTPf
4xuUQaWAH78dyr8jNMk50azH6thOhO4DgCM51Fpdm61nY8mSXdHlMUT9fgWKRCfUWUm+fxj3SdPT
aLH9QWOGo8ZdXbbkPDy714BoVsK3kxT5CDQeoBGdXcZKEhyhGVyh3gFcY9kSUM/ZKNPQXNqvUKQE
/viE1ND7EOEOJg1mNlPmCC8NxUVvgILbHakL1B3epDdyaGqMKEBgFflNA4BKZA8HC/kzR37opudA
rQu6J1kkARKPiu1iLydVPvz41CWUWTDZ8/FLd6cgb7i18lJ+XKmTY0hhnPAx7ISIS3pHAhAPcujm
VSLDTfNVjg/D4zwdvQCjEwKNVDzKZ2elLYyYMV2S2sriSG0q6aeEsr0+90fdUsCOPa+3isbGjKmi
RrXK7MqdGaYQ83QWWoeewoeK36dvgAAAmYp3n0UebPprSSE/1m5meLJ3YWnPgUQnjQ+leRhUsrUw
ooyMg+LCCOxr3vDyEberPrMETH66RmbxL6mLDTMfqRISh7N2/VjYnWKUvXlffgFTiJ1N0OAD6bpz
h1A2T6N542z6Q/e5Y+FyPw54yNGwgzwJL1JrxCUdFk1fCZe+HM56XdN3PxlMqiPwTHGs1W4vbWwN
TTmpdUN5Q+VqE0dkZokHyvOek4ssyCKqQOmRq7tDAEPwCZB91eYI2TPbqviDkYiJFyXYmDzJO4bz
fW10FE5Ag9o+gDzeJ+Yp/E9DrIfbHFrAGotmkbYLmDG4/6GzMZO2F6nkzEcAoZXCEYrq2/vdqHr8
FUBvA3ykRVdIerZfqwIbzLZsgPSCGVqjFQxHxC8qi7iPt7/zT6Mmcms3CylpKIIyIchH2EbFqfcQ
Mpc6VatMf5OSMV4lYku2wSVOrntBIs5Sz6ElL34QHkukgWq0DXWnrsAofg4cfdY4HaDcsmrcC2gS
M9M8pYYBRS+Wru9rKcbeCFHsNsDFADu6nLopoeUB5FYmTB/1BV6p0P2ji4OoG7j71LqlZl3kzlG3
oDQIEDjuth6i1JbhKoaWMuK+G2RGWXoc4+QH3oJGee2n7v7eExcPsqYvoyMJBUZRXDYVqp8zq3W5
MjSZxqLMmAgSAEKumd8phUqaWjgmzmdbYYMCg5krjdmenhGKTcWHb3y0pfQ4im1quDYURkHFC+1u
i4su56aLEPQZVQ9kcrorH1mXgO9WybKDZNvwNzPyO1WpuXk3+5d3o/Ra9N6/tb83/HMPfDTG59St
UoYP4D4KwWgeziu9Qv3j8ZbqaqR0Hokjf6ecfRemy2VaVOgfAJPH8622ya5C0iiYqXKptov7hzG5
DpmUkG1F3dyOtjFvfbmb7h9VfTVimY9XbIrlJ4vm0OFvw7KiuAVXShqKIuK2NRUixeR+kpM2ic45
gKVZiAL28YLx8HQUif1ulD28BJEgPm/M9nerhOjAKc90I0tQI0TqYaja2VP8DIZNy/gckhxhfOyI
opZJMReCHBM2QK1bo5CVe4nDaPDN/0WfxAB7LO2TJgUVR6SD3jySxxB+KIKiL6BDZIhBVnw951lZ
FyQXSSGFVkYXtX+5F4upsHT2knxAta6wDDaW05ga6RPpmc2cAQTpHR52AxT0UHOoxPZRi4He3XMB
nWf3erFj9d/HpL+nN7EIHt1tt7jcNVi5QdvW/6ZnqI3nqO8F26YrMPrwVKGXjBsr6Q+aCj90HGcf
THNpRs7G44/CYlzDA9zbNnqWfyBCmSuw1KtB9xI6dQlh4eythHvR35t0vNetHr0OoU6mk0jrVHZv
KQRNzlu9wKMsnvckKl9PWOM/tHb57G+TY72mM517nVjSj77bORk2BayTmLPD/SvRtjmkG6ZVQEc5
di70AU8LF4O+FYYKnXx5zbNoeXUsRXaAU6xGop9T14ALihq2+9UY2LyyQ4nzcVeXf7wat7aoJ7+Z
b7p4DQAU0JsK3FK9xlLfLPhYk9Wv5c3vzt8rThxaJKO2H2OzlM23EHv1BTgt239uH1EWa/zf+Nym
UDJ0/4jbyFr9wDvLJ+wxUPAr4vnQZoYNbLTD71x2SCznv+B1Lo2VkoB8JR4bbWqb7COB3Z3xu1rM
hVkLyS6mirez7iXYYr7xrQVmq6tTM5PGt7Mf4mI62fDUzQNOzLWZT3qVzj6tHViWDkRNq/MuqS+N
YA/VZbnSk4/C5c6QsZvAyY7gOuQOkYxRYrZZTAjCK2k7sb/B0EWQ2B/gYOnFScwm7bGG+cRgYJJQ
7oOpSnpgcGWr/bXc+WAWmhyB1ISEgfa3TpANeo1wGM0DvoUBEcifSuAkpTx5w4HOF5KuwPOb9r6a
L+gtf24RoACVzoOSeEK4A+OXZCxSJybrK7jwfE88RBBmLHM0C9wqbr6CQoKgIDUvxrX8uFQZxy+c
VqBNxotgVXg4Wi2m0o6SPoRIVY366ySOmfMTrSxx/4UK+43mKRPGxMiRmYLnDO0AXL8reNsgnV6G
lK19YQH6I6H8uYLayZ6Tf5QJNvdjkFvdbvZHEm0688YEi1P+52W8UFxoIezlSoi2U9o0raN1ZIua
co4zt9JyU74qFUCJogQtqsN5r6fMrypVGUVOQ2zxlyI0YMyV+QE+tmAeVtNc9yl/EoVuQb3JLRSM
z9KB8YckabN+fY7nuRr4qVlj2cBES49wN8oIsTkX8+G+UFSoLD5+Fc2UYgaf47v6+ga3q1XXngwL
0zIS43C5tIOFByv3E8/aVmSFsWwUrdqqlA3fs82hssaFz09droLaOA1eiawEa2VHZxepq9MTGGKv
s6GOBE8ORwXxgvYB4Arov4PyD70C1ilQIg/+cA5iLtcc6rIawI08lSJz8oPN8CcFRtlyxZnG0hm6
+tsiJfjDNSqqbj/eIg/ZGcsxga1kYDYg1yLoQcZNAKQWK0n9JSrf9KdH5b2yokZ/iBxsG4o+iFGB
gTxf7hu7JqGGuVb0CI26oGdeOGh0AhEz4S1EHpKQgmKvzDTVpPKexLzxtLmTt7A+kFs5Fl5bOYEb
kcSvCO7aeau1nXoxKeyhvOdTuldJ6+XAdhN4kL4OEuG2mx6chXEzI3a3x8Ww7OxK5M8ZFGu8kFpA
O3wByrWEl0u1uGKYRhz/9VXyuYghJilkIwarGhWVxi//8P8FUkdByecy8WTceAdOnKAibS8jAxhn
KSe2ApzS2L0NaYGAYzZdW4cNJWBP41frnj4dVBFIGT3Hy0z5VSbOF34lp+XBJ9v43ns7iP4IuBYD
1nTn9JFDxMWVV3TMQ9RyJQuDxGvDjBhCDy4QQ/EzpB+LWLQQvqagDNx5PUKilxx4mkz71oD5oMGQ
sOkhWwZIJciZBEKD2TiQwPc5Cpbf6Y2JK60yug6qybPtWgXooMlrt8y94PHgJknufSjdxrA0Uk1w
fpS5t9167Mb3MJRkzptmvYdcC7oc1uafnfh+l/bAB/oVXTjOVXZDfMDBgXbp+UqDtQ92BY9CK6hq
BYn18IrN+VD536B61f6qjuMfg3XHaDhhfnujRs10j4b3mbMQSHOfAuwHWrDZ3JCLtHWAkU+uRzXF
+Z8HsdZonmPGn5oFpexP2AJ/NangvXH8oTlBPtPI1hGK1wi7Egwjc3OrGuHQhQ+uDY9T4vBlTWE4
MKZd/pxMUd/UM9uXYBZgieot1DXKXRk+wgXrYAjFGUyfki6ek9+DzGrMwVbGKGoe97i7EZYHCx03
gmwibHVltHIlQAtg/BWhgwz/Yo9USixVT6Hv7nxuxki3EJFZx05xzvDpsmV3QgRHaAsdxK3ZwB9v
KTlsjFKZ7mLqmW7zAS9+owLGU7H+Y+gSj7ysHGHjAKrGV9k10iTZj3zHLDenN+1zbbg/YskWfja+
NIn3xY2xfUiGnjHWoOOkbipSx929hI/Kk+OlMvb3S6SPNGiQsn96RRCFLSMtrJg1nyZVZrjxRwaM
rmuToh1hM3I4NkjsB9S9cbW3IOWiL0guBx7P6RFnxpM38uymjCoNZAQbfxIHAVyfmNKpmL0V7qqU
VkmZmeLXWW5jOLmA+6nyWE7uDlt9VJL2Urg+oJ6wmyvYBK/jrInOpHDEWQcPCy+5Dn6jiKmvpgJD
akxUa7TVGrUPq7ijyWMWE8w+eXHgpyQp67sxdEnHtfe5qZ7Cg2LOTDUmJQPBcIC+YbWEk5M6z2JT
5sRICoe1YO32rTIzxTYXk3HEMGU3z7ohpFQn1UQkjs1bchTzwlBCr06UoRMtqMcmtA3ajK6cZGE3
2EJr/JOlUFmzdjPGri5Q75tgNxMhGgQoNwD/iSZTkch3165gfsVh5V/8aJofbyaF3r+UmF41RJAN
a/91ZfU6iX8TwTrDMJ47ukbxPH7waxQpPNXxHg217ejg/8LwYrpVrkp5aUBFMRr8vcLYNQkO63F0
3En6SokZEUxGWILtXHlfn2siJ4u4AhMOEwcoipEqCv+OmHxxqFjWBzzdAFxPcSqWTqn+2jghj1bb
/8rMhS7MVJVoXg91T5IUf2TFVNXpDy5xxElZwGmm2FYZlF1LSvmLMXQbbNgk7mMCf/eKtnvslb+f
uQBUTj+P364JIy/pmN3uUHxX46fAM1swSCmfVIUqEM9abJsjZ0rgf/VUvlVNHgA376PtEYn8M9Me
isxaSrUDYzX7RxDD5j5rekELmMCma0AaTIhThOTrfM4BqnfoszJ2ZNfDlcgTbCVfLN8in8HL8djQ
3IjS+JYuLbQWK/GI0yeenfivS6xxJK6dmpEuYDRWScEkkZK40hBgXDEOFynXZswNB06VinURSaAj
tsIhJsZsvYoXNxScNgSG7r9eGp2LpHdazoHweGxLilgPOXoQKemszZZGX3co2OiluBYbP8/FI9Vi
CqIDCLCNPRV94M7Wxf+7aULfvhRXOeboozBEPsGVibaKMyfoQX9Lo1x7sfpkpiF2RwedhC5Xym2d
kKKCV0XCik94OT5X+F68Gls+LfX9wPNOVbenN649ucggPW/TFem8XKMJEySRDQAoezP4+OHFId3Y
pPlZ8gP1yLdFL0sZJwORziUUQdkMwGWkyM0UV3Yc/zD+m3M/x5GPzydXVMRLz8ooBG+1r5wZSPo7
rKhzHttRvL+7b44MhpdkqRSS16/jRqLoTRIC+XFanfuRFBFJaGKdzDFvDrHLdnhTLiLCNd7u7kD8
UGc3mb2g6kBeutUPw6sheiFuOEQ5qVnQrPrVWtoCU+8EKxXMUaPsH8W08Gr+DL0MLWewZ/IK4RT+
6CzKA4rkmXjcauIT8gueCaiPmGee1VRmKQeE1TbyfsTIrELpZfj4UrCY6uVPUzQkyByCzKguBvwz
xsSZrImQmKFR9cVRU+KVYBNKYLHzEr++QQvrGEPpU47RjmK0ctClRS9SDb0Kzh8a1vjsPrkLuJy/
mkRvTQ0MKtoh50dpCwop4vh6/HK0llVXxg29pMWixggRg3se+++/C9aJy67MU/Q5iFh58U1yGVVA
3YKuQ7QFGAJhBzVbkIZQaF3ijb6gDQOsfbfEoNoPUXta3PWn16huMqvHvsPlDOMFzpUEv5NC1Js1
wfZUcTrzGm1HToyv7Zvez2gOKn1EP9ckoxh2tHiTGEG3LPdXwHdXWQZ+A+BwwoOViQggQ3JViX7F
bsfl76ZgUO8vGodK1m0m6W3IUhAv9u3vcvTsW8we2frGocl/pyqXfuikMfdTumlMIxtEvf/Isw4T
3/E25CdogDTwR4NpoDFd5USicmFkpAzWTTf+TFzubgBUhI6juJR/OAiKY94QmbWAwDMsVkKd36YE
x7jRHWdsp85xp782y9foX4F4apOUETTm4sjifGuD55prTSrTKfP4Fw9fFG+Y0p8eL1fKQgL0Amqp
JLW5hcuX7vtiWBSLFKR9GM/9ShjUTtplRHzSY7sMBfalhNGkZH54LYbj2d3etAKvp+jZW9XBi358
jzH1kBducgf1NbM6P4zmdAezBtVEj+ePTN8L4/UwObHZyMt9RwG2Ytk0MS9ZggWXQ++qJiWUvV+J
pDATCGhxV5yTbmDyxC/2N/SD3TsFwivAENt9DoOGBodKJL6uIvfrOnJCaLeQvPFdVk/Za+nSuM1M
PJZSYbIJLjB4qatN6xLW3aOQUEKDPx5raT2FNsKOhNI7mU3gSuCMP+F5LLV3GHI9nE1kEmugFbcq
wMUurpCkV3bdMA+doVyzqUwv16RxesatfP91a3VMHYtNb3ODxc3tW+mE9VbIwWeYIM+IhbYmvJW9
pidKHd9DNwAHR89sFjGk8healixnUnjnctIqYVXFojN8/bNen+tWEDmbbdx13rCXisLHazJcX5mV
jsim1YFPM136Vi4sdI/+3SQQICTUrEffIAtx7EcrR5h6o918mYEw/SJP+ZHyG/rMWGPp0sgNRREB
gXLtaiHr6HJ++NAzq/s8v7MCbOmBdIe4uW3wpIHXwi+vZlIRRwRsdU9a7ron2Hb55dK0yHnHNuZv
YT6KCr6Tbd/0j8QuKJ/jmAWDWTPbUV2fbYqqTTPyRi+/70HZ2pT/XM90HmXVgOUfDpkFgXmeXEcD
VQC8ADgmfRSyQ3M9ha7QQTnL5hApO/nLOBejoMMSD3OQCgQ5H2W1AbgsZeHBbmCIE7X4ke3SB7bm
/Ycsz+WlM9C9XP9o5EqmBwvj07UfRk8yiyMg/DBM/JGOI/rocej99GHDiDrnW9JntOhY1TV+snEV
lXA1GRMQ262R2wDVnM1FLkUJYVFZ1WsFRGnc/w9uLXL7i+O15VguSesupDbTkMttOo2u+mo5a6s9
2gitFE0k3rv1fLeukgSGZcehtNfsnyHQd4DAWfZ3w4EJxTVh/iBm8b/pB+8C3Br8vYrCO+LZO0Dp
0I6fTe+lS3oTf1HXqW2RQwmI73oe4gXb+7IWQCAivL6NdRRs322I9npZHbOOYLaN3Q58yC7B4j09
j6AA3r/TzPuvN5giMM2V9Go7fLauScEuqOn312Xo9TYv4RcuyvFHqjVm76yMJL9TVA3uSvXOE9GF
RIeenxEIs5I2Fkvxvfki19w6PGtDO2GCj8QZFIALV3BAiEH6x/apDjicJbwfbkp/3wozuSlXbKHV
n1R/ZkYegTjoNRfBInjUOK2uLJ2BIezk++JRXTs4Ci+sk1pknw6NlmoQUmdNyuSKzXhSlzMxWlb6
7RMbVKVmFyD/794b8LHRFJq9UewrA65V7ONrg9uQmQQpGSk3yF4bJbTual6nrYgyBC/LpTBpr6Ma
55GKeWxPKnscGY1pWKiPfDqwZETF/uMIV3FEjxLkZnuwLDMEUX6fPm4WOWYaI5I2LWyMCC+RULTB
7FyKnLSNQomXcBGeEUXvuz112cTr86sS0si3zKgXp/kcdLcJ26Gz/JjXZfEZF5B/Xadokr6N9wQ1
GHiRujLwQNzNNhoMqSPg99YyKhL9SOyvbmBmuOmn0yM+DSOIRxBGqxTgA7BgcL+8J9CoLIec3dVd
FgjiF2K4/shqjah+k1mmE0jUpvjxOMCbBEytHdEy1aBLAoqSaJ7hGJEczQjSu3WwJtikVqBBhWvO
4Ah9z8esHe59YaEKarYfMWIopToqIPjijl+CeyRluDZLBfgCNLwQHvpMUfvpyaciKnfkQBAHLAhI
XPO/9rT/N7D7R5KuqGzwqKIkXrO8wxZMn12G4rwRQuyxJzoffONqS5omM/ExJ4GxkR4G5s2lkWWX
IE1tZFEaQZkzyvb8jiE996on0hnrVbdrWjNOGRK5SrIPH5Q2rUa9lGh/xIJ4qGdMi80juRr6ZyGD
jO2xmD//BU5cZS1x7fhrv62yrUuaiaTUDDV+um5pm+B/f+KiDOPShUrUs1waDY0cKBm0q8YyA0HJ
K7rLuL4lg5qvfXX3qVjsTHns3Jqaq/spfsvlVAZ7A/AOYuEx2t5R4QO6kbtWoh1ud8uXcpWFtjPV
MDF1yfkwIGfRH1DBeU9rbPfIbl6TgaBpbE0dRc9iS03LSxbZ6Xi+3kYX/AU2NKSlgYZQazBHlQY8
45RJEABe+ME0YfdGcCijFOfe38XxgSJ7zEiVT7iiIiBsdctuhkByKTUumefbIBFFUGqQhKvKh9Po
G4CaxEjmDIB2o3hVa2hpNg1F0bUpunPIvmUMwV8g6PdfVnw9207R97C7T0DZYgPluYauWXV3SzoM
LSEKOHnmXGCVFHYMuEBkn+VaEalPDW9rcpWvTHcPzsmKW1NP0ObFRlZGiX0foTg8l4qQjyjmq+fN
3Oe01T0SNDSOZY0SDRlevsY4ISpjDmwCdeijbljtoAXTjvko9GKTm8ZkHhswZY7Aog5t4p+gdUkB
hl3VdQu5a+cAJFXL2k21g36Rj/FuELLGzksCZ0KKgJExcA+bu9EukaQfp3Hm5GE0DKRmaxYEqM4+
O4LzxOXYQKEtQ4QlntbVf6XKM8bCIq5qdDdP7NKrQi+khkpiHPRt9Rm4ihq8O+hn01Nw+b58NUUC
GFTqYtzHgxV+dX9J3z5nWavCV9u/FEMkzobv1Gdil8P6CWkqvB+IZLRFkRJIaHxloWLegXFnu+wO
yGSylkUEiWVyIV5Rl3/jFJHE+PKbIWaz1/0u990OM/tl14lzQj6BjuYzr7MwsIC73xScDTEZ51+R
1JtfM2s9a4TEPbBTK6TTZxuAhgdKvNEFTXJQrX8C//4l7cVPzHR75tSg5wKQm0Q/1Z7s6h+RNfCU
H/YtOfB5z1yJjFINRLeTVl4vyD290ExPsBGYpQCLgK8rNimbj0ok2/06vHiU4tFYT1x7JZ2vVww7
EOI5r/H1g3VrwEHGWMa5AHDHlA421ezOIKlRR97niJjAHTtMMC5w1T+QIjJVQKwt6UjECFo27weG
SAWv9QcAHfGsTTyzLL5lN0X7Ne1jErCezl0mL0vAPhVti48aLAJP8P5KWbkNm/rYtWo0gLT/pnUE
TLV3JX16eoibQSAhXpStF6PxITHXWT/fZ++a6gyZFVNxuTjNy46FjCMSlLaVoGSMaDvKEE/GEtRI
pBAHwl7FdruRpgEC1+vjZaaJx1LDo54RV1phyJP+b0ef4fhxflhySD3+evbGzidbZo+KB4oWTSG1
xJKlre9mPE9ul2UlM66qMUPGLMEvQd4at4jSzzcvesW4AIgw9r9zlSacH+xAtEOdr9NKa3SBCt5I
wcgj3b1fGkdFh4DYjBfctKBzfx9ByjxKPn9/blscfniiSb6O1nzHoZxKcxiRme+VG4YV65NYX4oq
Jzq6f6Jvj8RLsLuEbLq2U9XJU66S5d1ZJvuCbjtzg6n1bUmBG9FcdNry2/0RjbxlYH/KkjYHjQvG
j/hE9yK2wUEVjNHbwYE6n3Q9ekuIhoXIVGoAe7Pgk86ps3IdYUTxXLpFll1QZYOx/cRSdI4I/IGS
KwsVX9p3oJt7EP5Vm6p9yLeIT3NoZe/w3SPG3UJ4KO6NY8NuGWpsvIE/WXT6LISriDQQTKukI9Bd
zT6HwtaOK831G6hjY7H0IhHw6zB1mFG3/yguuadAMrcg+o2FCB2u1DmPVwciTtaeRa8krfQUpBGM
1ch4rqF4cv4GQZmOnvGd9gCYBgrM33nTL2If0iKpjltollbSM+OQSZNYOk42LBpNEOYDGQ4YQr05
0js/mwW0FKHrL8+XvU46bcZXMGJqJDPqYngxAa8jAOm1/ore+W9s7h26jJM7fl68qj7P+HuejoM4
TijRZU7u5Q9TBrjZVBblVHaVpgUGNauLrWc8vgBOp+a6+5GXPV53OUo25kslzTEy64oYMuWTV2CA
5uMIHeSSFK5GmC+F+WloH4gXdWzDKLZWWL6bNzJH3uyIoc7Udoa/xBB3Ylfoeipu7Y+jUhyUCbxe
YaoWIu//DsYkTDDy+JcQGM407kuji03zWOrGFAtevboR6aGLv2uUr4XnbEhR0KA9wE005j3uoqHc
UWgEAygy36MsZpMMFIMgKWa64xwtyaPLEuiHZavp7bg1KNaAoxwonAsl0DxevhPR0Jdm9pBOm7ff
fEocYS7jw/6puEbNHvc/1Fgk+P2TvyWUtjtFvAGBCNS2/gdI1pEScTQ/Yszuja38NMbPfA/M6VeE
5t84dAjWH405ifj2cSpnGZbD8ikYivRGbZMTp0jxTAkqQcim11DI9zCQ9uyn6bqB54yxYATGLj1V
8c8Xf86LBybwmcwXW1Ia62p8YTNbiqR1zTb5T3ea0OlA5feHvkC8KgImcBgvrcbt+Wl6u36qXC1k
Pk5dyT22g2dxnZRi7rWeKvcuJ9feXr0VU2H/9jiCwEe9iulC1GnSdgdvK3KI6T8sEjJGuwJHR+Q3
W9jrajIj2T2if4yvuQsORBRH+q9aw0zn4bTJlfWKlMSX/BOjfF7Lh/A0G1zV2KzNG9ti1SSORabF
AMqMY5INm12VEkvj2o5pD0i3W9LcdS3bgJP79otLLIMd9v+OWEciVKFNrDo4p1iJxVTh9eo7bZYA
O2DzkXdYDbLJpLoWN6Jyg0hi2inPYJvsq6dqXkzp0Req1JJCrBVC4+MONBKsC/zP6gFVQl4ReC+P
DmP3uJRd0yKoOHse2Hy/DGgKnial1m0gerqmVEtoF/awEUI1ZTnMZLnRkOLy1tPIPCZEs4rq0JgE
yMexPGxBgMxh6xnQ70Zp1RwpAvJwdKSYL6CH9Gk+0C+ldnrxSDkWibQiUEpOgo7oqeBeFb6MMFh5
V0wW4kGjk14IInNBe0GlHPHBqPCufn9/mONjriUjj7xxMznvaK/5o7wRCz52HMlXKoLlmULrdWj8
znSQogFNCioB6TVqcXYMRY2U7NbFutEhAdfsnys1IMhqqULcxzhiaE1+Xi3BF4UNXv+RmEjUhc98
U4BH9Xfn5gr6/UZWgFMvJO7uSpt5b7XbaxymqiTYNC2Z5Xue6/3oFK6v5tex9onztASIsQnsGn6t
7yG+fkcPvN6DTZMwGElsoLPPZYsMW8n+XlrWgdfNnRiHj/viLsSlTIoZ6ZssieWH3kzxGXSyjsW/
lWaaVVSEOor7H1qYe8API53w2aAfBNl9NeH+/IuPb0nQIFLpoj57XflGdVwHm6uEU327e1QIZA2y
3rLBWbbWSGTa4EJqBcBGUswNCLT299MwjoxHVkPf98DcEBb0BJd14CO8Z9Fus7dWIx7BsV8hUtDC
fPOG3u+/ECzchKEbcRmyIYidE3MREnQ41KRsgBGnqohOQKgi33Whc4Qt6ld8OCMHO+KQHaD92HxC
0a+242il8HAoPjJuaWYMnVr8p/2zZwISSnO3rU4+wpmDKdimmqqs70ot6sPimYG2IPUSpBjcB1bl
XhUpUyxHaUuidFWH5A6g8lnHTXPJlLQwpiFrJ9uWTm49hmJgAVfBruKDBZQeYWy8YiQliQ7qU12a
kvhUrmD3DnCl7210/gxAvgWZOVXaEDzYld+5VgPce9P7VA8hmmzOgzjRbF4VWu3hxbBBRj6lThYX
57wbpgqv7MuAyq9coh0wOEgJzU3ZkJA2ZCeBEey31VEje1Zsskcp9vAhKZ8C71wnV2njrAp/+fk/
OTwebOUHfJnNxkeYps8RI+0AqbHPNbMe/5OCkXVV6DaXXGy1fk4o8JFcR9dGhWKh1VjKFwigUrCv
8ZmqZob6/7bqe+F7tIakpwPe7LyWgwDZAE1YVx7LMlfFDrneP0WaLuQmuo5wzGxh+9CcAdLi7gR4
j6h6lysgPp6lrDUZa/vgRPy8nP0gWWR1Q2cxyG/MUPs1Epa+B7KDHDY6n66XE1TCXIaUHAQ7Q/KN
fNLEmb9UIN0wc6xqLHJXRxCWJqBD3Y5zrxqIhDtkysnsvdX4rawZkqwo4NwuOgHhTL/+q5CLCNJ8
XbSDKRvOATltKcpC2/DYxh7DqjTOwh821xqmxuijI3ynhv+sr9ToxmqZBhpt86OwvMG+3HG+Mk1V
3korfDT9kFFuZ4eyM6Z1uxvLftOZZAfVQP/zft9jmpW58Ldvn3g7tvpEB+JW3jbgWP636s0bxVHI
Y8UlYN3p/vlWx97zHtPTMZc3OysvgFsdGw0ByhzYb8K+pwCk+tj5vhVKsohnjzsDSLWL0lQ+XPdS
PKcMI92b3HmFfkaI3Zkxiv5952cH4f7vbQzHlubcGY8zpdFSEQpL9d/ClRld+9BhHRUkfUP7W2p4
sp2aBNaFPXCmFi8+XChJ6XUYrYgGegHqPawiSe9LVGZwBHPSCtTcnpK3XEeGQR3/rCIhd3yLyT55
zoDoglzWj4NmlvI2iIR0M1qHAXsl/y1qNHvcZ2/728KdFa85kBG/oo1WZLQd+2xKOA17dkaiZytX
ExlAqOmqxUGA9VL/BrnGP1HpYBKmkDwWWap7/sQjwUiV8PN8Y6uNQmA7eQNjHJEJEcWvBkKDGDB/
z5tL/bm/n1Qv3r9/A/Dce86aO6LMwubDYKu15/+7426tAiu60ulwRW9vHvv0XNgG77YROaDGd0KG
U0n2iXV1M5aiABXtv94x70WZY9vr8ZjHPudEwpEyt9/4os7jdKgeJipJQ5i0p6N814zbr6SO3I8X
Ll+5K8qGgsziMlY+ujyWPujVA938M4PPzpskaWP7aWtQHLBVoHE3jq1GDXa4SeSUfsgWRZsBg4/+
4/8VE+Qe6gnmbKIXArihAe7h2yRYobRwXFDhKy54TPPMxdLfjSLaopbYujd3fwJcwt2xV410uPx/
e+X58za8XZX1K+pYrf3rlFDyTMASlz44S/2Jm/zsQoVk65NnQHXUmQ80W/x0+kibKRTRF+kBPfCV
Th2utJ24eiHKDtUK2W+o6zNCLxe1Vhvd3nQ/DuJgQvijjt9xREWb88yu7CkRL2f5dT3/z4bg+alc
8qWJGpfdJeRR0GFRHbUTcMQl0twh5nnExJE7+GIHv7ydhYnK9C4wGE28RS0qVMzSQi13uykFJ9XU
TSVseSFV9MMXhVM25RaWsR4p2DV+bSX+5pv16g6KZsfKsMxiFGDKBVCu2IAZ8afsIv6sD+pkXha/
fUoMo/KAeFpa6Bi/oKdd1t2njffdS89HUw5XqibqQ83gWsRAEhVCL3sBgwAZfmJJom/jgtuGw5OQ
+b5H6gVkNESaprqmAAlJ/AgYkvOZWEc/H6LMiO2mMQx+0KMDgXh/v9HukGt7l6oC60uA8G5bwyH7
d9IhheBmWM279gUCNalZU4Puufe0ekCRU4LAJw650iB5efmVpn+dG2QrIGGPI1waLQlzImGpHqGL
RTH1XKLvGV8+igYonVqFYi8ZJUNSbICX/yCzPc8LSoqNbQ51IplujQRDpeESm7y9qu1zLTelWLCI
BgsIQrJxgEAswR9TJd/cPyoMsLbaP4T5XvlCIHViB9ZWv+wWj/dTO6BzH3iQMvuH+0yGI8IVPyVX
TfPyF4t2YMBbvqvzxVdXlrxy50L9jfzgw6VorFWNnLcX4c8rjhCNEsKkGF6ZdnFGAmopp6pNostB
ZwKpy9L4YufVawX+mdKDNCfmcmCrlDSya9nlM2dyq8LfhSdftxbqWy5q1J8/R+h1ep66xNnYSH7E
5iBFKHMccFz/sqndpzzrPNurIv078CUAcrjD9YqyihvYq9JFpntZtJh4WBDb9bD8eZHn9v3Qx6tB
Cy14L1FcHdOvdh4mv4kvNj/PvGud3ddv35pnbOHeaI/I+KqhnKYLoc2XCfyjFkqMDGTifz+736JB
0ZMqYnS+xP9XQXdfQZfb6PEW6yoChF0JKMRAYRTfZiQhZx3Se35ypu+HgwV574W6fRxngjIMB7q3
jvTmp1eGKV6WJsH8bWMTLlS2nt9H2VTc026+e0KyuyKAEVK6Vfx2Ry+XvF56HUPbQ1Jw0B6qWpb1
yDtRInZNjiatDC8eEQxXqQrA/Khpc0D3HaZ/Y9F/a0RguTXxUYrZ+0zRRJOiHbugg2XdSRP1pLXF
GoRrDU2wVFjtI6jtncoxLfjX6l/jbNHKsVpilFBRIEuJjlWgCwft4PH4mvdXn5cpX4AairzryrCC
1xD53rA3JFTyisnUPQ6c12iHrJix8W5tAnl9n/BJQ95xztAyp3ZjK7hKaRk6vxPvvW2bAOOSPWaj
BV+zjv9J1aVshV8l9thIM0P/IJb9a6LZW2rAU/56X4x11uKvRAWfENSWf6Ir9weZDfnQYSSzXTTM
M1hd3i41Gn+lrY3HWHxQuFe4+7py0168reKoiDKwsDe6OhKudpEs5Nm2heGqbHpQP25ufCYn2PAN
BAOji7N4phLwA1LTb2mhk90cex4zoSABGDMzzA2aNvRwWhkJtH8xauPhfq8P0bdjbqMpR5m3qQsu
anBeJrmU5J3a7vpNYubSX1CTTmdV5p4aLF5+9hKnFPHqvkq8zjY2q3dp019X/RuP5ylWq4Uo+gRF
5QLiDu3MOxeK9jseZxtdfvIfKIjbtV/1MaSz5MwfkPAbMfCjZcHxzMken+qgcPNRBea2eyLIfKvD
Q/Iq5HvyAoHW6DxSOux+crIBe2q3QEoKv7+lbye6GMQpDU/PhHeRODjRdXzfDTx8JJAJOQs7woda
Ewr/7khTiqF5k/CQCMAo+Ybmv0wyQWvUae3H6NSvlyHkHd2r/Z025nTiS5u4AwMQ5TTPlPSOvolB
YYfqavobhomNMUe9J5LhVYiwxw8x/PCkBSPcEyOKVbpZ5T47R2/ZE55lfx6gcoy52DUBJHriQ+dt
lL7Ogdh6A6JqYEohVwrLsDAtINjeKmHvXGI7TJcOYXDKYZmWUw103VDT5QSwbWJFBB9oYYChS/a0
72ypMXeCIyYH9bnrXX3OBLSt96OTecNC7C7SraNKpO4XTkj/58mNa/AT4+yhbbt/YO8yfgqYHxmS
a0Lpu2nYOti/oqT4zurRiBtT/3Jp5ZiZBCRZu4O2SMV+f12bR2dakZsUO4E+h4fjPRUugihC8G+0
94ap7T8w/8xtJKmRUrQSiCoyVTBEGRcPLZ20B2MT36ECYguCaPjA14LloXLZFrNhcE0COWFTG/hX
XnSKSxVoGzHH3/toKKwqUwjvddQ+FXILmmvUVg9lUHwjGNHMRl04Cco2JCUM91pobZePWpXdLbkL
mHBUCsG1puCGFRuKlz3H6vsqxvf92Elw1PLZ1/yJbBBNCZx7tw8XpMFk8GWc8kJXqPHN6g/Nhhbf
Z8Gp3qSICq3dczjlm+SE4bRE26AfykMD10+RlM8E4iESaGOUkwlJ9RTHQzRh6ok6+J4nP8tFxNSE
XnUhmrPxv2KGQyyEEG0g6/tcqeqaL6tmjA2vVUM/CyfuDBSo87ymoxGFdXRPA4UFB8mJhQE5Edxe
bAOOm3Y4MWVSRy/rT7IwuxXv3hrROdVSoqBQ/hgfvu7NW+j8DlbWKTXSyvODNXI5g0CEAr/F3Bij
BFrCKtujbq3QXri5AFLWcADluvgxNcDir1WdoOG5KyPS24+QQ4FqghZITHf1q+vV7+UlKIkJucZ/
chiPITxJtRod2fD+JzjLBwRJ6k/YVciHtmBkuG8cT4Q5aKocN25K2RBeZsyyyIqd7xY9VGjTRrvN
0YGVMxmyFBeqjSwtQBZjsXsvmmDh5WhaCUQDc//P1F9Zs9bCu74IbHtGlwLrnCql28CK6MclGh1/
ooJBTMan5dDUvztVeJ71aUW+wRcfrFTLsdLRdDwq/OyrQJkyQWL4Mnyjv3wpbXZAMKBvifYzgch9
VzEtUSfyvyVlYKe/ivo2/JFITC+15NiwqK68uXrUzI/dErlxwFj0pyDN2CvbLK+q8G1w18Ng5Itf
mliD0ixKDPFOBlquYoiZuA4akCWEqr7ruASxWVaKkZsWkrwU2PU8KlZLG2sOoJET8VZaNMe+5OK7
mfyZhK2lLrg8C2U2wj+RPsSGM/sLydeiW1QpStACT6bNFSbKp3z9npCmIVIrBOhhmyt3xPe+aoDA
TaplzUWC8qd/ozBH8PujSTosR8jM9Fywhj9Yo/aUcD3CK0o52XGQ+0emurRJGtOkxq4N+6aSh9nB
XQ70IZMpce6qEkqINHj71aG70jEi/RdEuxwq/17Er8Oa2Yx/HnnzZauTA8qhzvrqBSSeAcnz5+Jw
Gl8yH83xuBjNbtWcn6MLcJHpfnnYEUau5TWG4preIcx+g9VOJ3kqWLl/jTV7utdOHsEdPmuHqc+/
inaF4WXXTd3re7v0hZt+72p24RPIVGSXgCkS/iUxX4wMzcCafObhlQHv/LzZHhbeD9W4e6+umVJP
p/gBpke6C9xnXAFJhMN0M9TzCIGY7AoFGzChJ/VXFU14Hegn/TCH51aduWJInNtkf0jstcZYzynf
j1BkiZ9LC+eQqIx2dzsxC2iD68ncVfccB+qYgrBxf2CrZbBUtRXAgMmgc3cDVInNA08KBKbgP2Gk
EVNJk2VAiS1synuw3uIF+gSQBJpLE9fKb4htqY8wgubYK5gT4dSEfHrM0qB7kxGY11Yu5uBh7pYV
Lhroe3LXCLK+TeYp+g1lhTyQoyJmoI/kQomB2I02iS2fzSAen5HvdwXhigXx9xXqnPJLbmPG8Lvu
qwU5gxStkAHrNI4FOHwNWEVgj4QjLW2IkCV/WyF0cRAh6E15UlJvNFF1yfUFtMBqbSeH1+ab4vwH
CSjka2SfEklDVNF4hj1ZDW3+pAO5rFmvtzq7p8KpFcMZ1Iw2NV3R3SQTEA1B6SqBIxge64e5nOXT
/y5TGpyaU2D4yqHC8pVw78ZqQSigcVM25TYk7//wEGwOXqHUvP8iR+SKgD3jSLQfpsb/1OF6LSxw
izdQ420uW2GuJDglHJlfJ0Zn4vIEGTeWGxFEaH7rTb0SCYYShUtV+HrWMjyADyWeuTACnq9vUImM
d9l1goJcVxjfEceM8jB09FTgumg408/NE+lYf3Y690DMOtSbf8xvQQ+HV8smEjpT3IN+ELw3Mb5d
rl1y/oD/u9Gxygi1cds3W9TQiE93fuy3DUkBtIohfsvaIh58IhkhbnVYzhb6xoMLLBcaCakibpxV
1KFX9CA6zUiZ19DTl82j/KWuJE+vgKkOrpAtP0Zbriva9C2coPWM2yMn00bIZYtPzUuwU57EMNC/
dKOLPATjkQu5jOkuJ0DpxYMb005FtixUWTTpgQHHveSQ6ufUhixWZdRSTJZEPTBGEDKd4Z4u0rT8
kZlUL91dZV6ma2qWdvlb347uZ9P4T2QOnZGCXFffdSy7vg5st5IkyMlopyx2Gqd4kOM3feqJoZdg
/gAdZoWcYDvP7TMd3UiEvswmLeH2OAVYfdYSrpSbUikZzPJuZGRlaCrM3HPd1g+S9B1LsU0M5Ts0
B0RDp+2jqSaiWWPZ3ElOLsZdIN1n05y1RiTGBpiXPZzVLwq+lCflHuf46hK65YG5R4l35g3Oud3n
dIYV5d5ZuG94yEjMReKxZmNowfXU5NoFClgv7GtTUXPG9qqm2qKtgS/+OUB/Ux/RKD5iIno4FMjO
z3vLcHpfaG2mUpKM0QoopELZO2EBOrmLhRF745XDx8cxad1dEskFzkodWoksnkRdgh2PZwtrRqIu
2TIuh8QghmGbjrCtikWNTru01OMG9hb2O7x1ddATQ/wvSQc6CQZxw+znExYw/2k75XJRNPUnJlaK
Gb2RWScaJtZXeC+kSXDAhNqaD/dnPM08rFmJ+eRGTvajkJUAKrmRhhkYBtjwBq7VU4vR/44KzU71
fRpwsHPRicTPUiYR6CNBOj5YUmRgG218n7w86EWts2ZUnC19/iAA72ejOgACy8IRcySRV7louvet
jhEpKRegCvrB9X+yYbXEFrl20m2HMEBghG4betpUuYPIKuS5/fHTWIbSa/VBvYnLheksh50LYRzJ
9KC3EDHLPyHTXnJ9+JAM61uuSbA6iM9K3Kx2wS6XgkjYno8wKwiju1cF/WZPhEQtScxHrXndY9qk
BP18fo7Z8ODx+wWHYcu3hGDctfya+hqvvCu90ELIct1X3ykrIcA/jaNkK5eFghQDV0fU/XsFoceE
FpTc3mYPT+JCN6a5R3aFAKNy6H/WDtMAQmGMLDjYc5psO3iRmO7/Sl1WyCxqt6b0BNfcxDywl4/N
vQGfpW5GVFai8JgO7TjQaZpctluk2u4LSsHJ1UuiFKNt3p0OGHv8+rjbBWH5vv7WFbjomzQmmi4+
sKuaNCtEGQ2uHDhW6PBp7d5aj0EDpVYdl56wmmj9kG3Bf1H24I/ztCmBgSBhmGDyXojHWGpGLQ00
G5jeVUc863G/aw9NosnK/FqYIT65/QmadgBI3tAJlDgRRX3HJ1+mR+uf198FTM5PS6HbDdzF3U8P
QHgaJnyZR/+Oda0jRNNuQHQCAv0a8yDw63RCot5AYfnvSQxwty4qJhIj3I4WUYtv8tsS7LyvI2Lp
HTW79tNf5B7adTRBimwDVUV5fp84qjN+GPfLeAfdHSSUp4GxaABUV80+N/dYRNt2di+TZwHockde
wLOIJFeFD9F7BpzVnj2aKVm6qPM+TlNL6qGFginKVPPiBEkxcIvtxncg6uHBDf1WlaVoijySZNj9
rA7a5E9GAYhDisyV9uaXDd/93JX7Atx4AidDwGaIcpMqs2SYE3MH6ZYRMJOxwbvRr1JeVHv2aaVU
QP7NirILC9+4w1+YGF00Cwq9iyUNh9/94GBMrLSv86Oc8hBF+gY4yeP+LiXB3kxaL3/Km8gDg2In
RJCW0xtZofMxDHaod19liMPPdMb2iQVtDvTUzE2jplICyDzDnysivPgXOjUh+TlJIXa47lZgEObi
cLLTb6ZZqbfk5Yg89VUdlu5o3LpASeQ97Zfil+whPz6Hw0dIe0f7L3WTNgCgEv3Gx109aba45g+4
IesGRKq993aSg5/BXk+OQpJ2uIA6ngvrO5ebqkRleu1MoXyoRHm2y9l8pgJhisGU6PY1HtRj7D1a
fLTscvGR2LJSvw/JPMsjEaYg3bMDqqphy55cQANW0FSglP8ebzKRDrBHqOsUpkVr+HawSCuFj+4f
VaRTqbVolKiErq623Q30zGi70h7nfdI4WPG4Sat3G8rpqdWcke2sOhT3UyCQo0BSyrsCVJiprmgK
eOZsy6lDYxCFhSbjCxGgVMNC8YtiBRdKr8AKIZ6KkRr68SpOZNmtf+Awq4sc6kPMdxeJM7Sox0+z
eVnFnp/UxvcWE7rDI9iKIZDuRPRfe/cB0bG6/MHy22FtXFSNHJ8c62g9fCGy0HY1DwZFwKD4AJKD
QoyVOKA4ApC64OhsnNPTpvpeeLIqKcicQ8lrCEBmCTuKoNaJk4fessv8WE7wfthxNr19j+BueobE
KQPBegTrAuIt4jIItJv7rHDH19Dwmv6GZqvZb7/yM04qzZOJUX2jRO3ruOc0hwKE/K0/ik1feD8S
UEj4zecLn7AfKUZ/6c28ZWgEopKFilc/T856rDQ7Zw5JVv6DNOdLPcesgtEX7KC1ZKzNdWT/gto4
DhRL9nKrcWIe7eI8gX31a/CUJ8DTZSNKuAPGmNRKtfk5WPHnkRUzBQ4L0+wDt4Ne26k76mt8jHX4
tfn+Q2uCdHz94iZFnEsBYwUMmvwDguJVrvPowMSi0NMpHGIy0Ws+Xq0AMiyKBXnu+tdwaBC/2XNz
q92kZ+PsWTbIh+98iRFH2Zzc+pEL1MulJi/G1VzhSMLoJI8cUslhyIBesuO/ExeRysR+njGqU4e3
derw14FBe+wRSYhnbm1UwUOnkWMf/LnhsQe16/3h5d5x360UAieXla2IL+tPMvg4pfE4+JyC10bD
idA1oivMh1CKK0LxhaokTPcvZO1tSPRIZpQAqkw3jzMb7O7U6y+tIL7tYF32Scraqg7iyLXNCrdt
/qVUmPSVvidQvSNFdJ2w+SvMCpwd5YDdiC5gwBcBie/QNCHiu+mLxUTL3YTlmen0iMPN9+clkRU5
3HO60jrP6jgUhtzrpfdtoQ7985s9qQJasYydWK1M5NTYUSQP48mhZ/7XTJsEpZKWKbqvKXnQwATJ
TH2G5WxmN8zQkVOy8QO1JP8P1vQMPYXUO8VUaGbhaQJ14iJDRKXStrCAzPpb7tCp9Bb0WlznvhqG
cCuYanMxzdVsknitkiokotkSXVoEnbVjNGB7/O5lGvd3c1WRiRDCBc/0HP+NlFzLNnyCicBYJzmY
eNJ0itz1kubF4hK4W2B5XgSYFizHtxs0qB/iGDRoMiFf8DbMnyEniSTn21WnLu0l9SWVB1al8jHK
zIuCLNBvI/E7UOUdo9s8AoQbgQOxqaBqDoYYI4rO2gtTVRgUH/HOHZ4D097pUwoH6RwNdcj79meq
XP6R6czxHvc2a0LOC3Xs9H8w40QMUJlNKzoRGcBXzFY3nN0IIyxXqm5UGVqWhpCuksAuHjn6D6XD
lWsYeEMfsmx+1s4Jf1zfqyUmdW82Kbq6rpXPt6CqqrptCU8H/va3vGSca4dmDyAew/Z6Qm1l7Nzz
SdRXOFZelE8yYMv/riS4KDA8d3EfybDGW0Thn05nEsxu0owLsCzQjzuxbbFCV1scMvBaj+wNttF9
P9VF9/66BoU+l0OYoBbudQChBLEkr9iXfjgQVNq2p1zN6slYjODXa9vFyeycvVwqLhq9kSksuouv
cYQh8yc28rksk9tMOwnLSXkzTcHh3R+R/95JWkOkbsccCDo869WwZRYLhezObCstZOR7/2jYrUvU
RNZW2ryAr/T/0DAIA+I4LgN8KxQoMNGZGsMKljZ0AXZ5H8jEet0DfY/3SAHKWNtlLMjCp/ORMHH5
E+CYK8PGGa7B/0WHm/Z+lqxuI3aKRTGcOIe58uCvNogyL1x9UFhDPEV0RdqW2R63Nc9BIaY8ru+Z
v9BjEGxm+mCkwPGRoITr/FZpDvmJp4IIvS/g34cm0sK2bLP/35Ug7b8o5OzeJlJfIY9c6a/YPj9j
vyw0gfRyXQtODcMgLFK+pNGOL3p365L1YYjKfAZZ/uxZF0XRZJjUfAWFFKR+GWnW64FWTMH9lTZ7
3T2wqS+xAQ918pBNQGzbHkJJs8YAHCfG7m9YQTzroXH8Ws0JMzmDw6NJiN2tY9wNffjXJIrrlGuK
2SdodMyjDbKaOShF7V1DkIGq4+a8ODe9HOd+dy7eNrfMm9r+XFNyrL7he0OWo6Q3KFKm0Wte9DSr
1q7CZD3jUu+cZuCNrpPDXxIURD1MpPtJr5voabttwa8E8rpQF/9RKeCOlLb7uthvof4zzwzIK+Nk
yzDx3BpgV5ZgANxIc6mJW24XT860f3RN2cQQs+fdi8ukT6KaoT7MvNTAkw/zj970wdUeYfrZ4x1B
Aa5gTN6SZWxEMvzqImgyd56SluFHPtpcspWUfpIkQMSTZoabOOYRW/MJ75j4N8aDmAflOEGjKczP
1cuvdOPgHth9fQyPW3y2JVIPFiryN47bKmhrSxz6B5oM1mWdqBwqyy/dIegkhL1CnKa8U2WmVJpT
4GwlVHARuoMeYGXA/RdHGe624beGLl4zSojTcgs5Gwqn/2ATEuCsqUy32TFJ5QwZPZPvpdb4i2oF
CUTYSuq2oNfWhcHsMbjqRzumV3zZl5pk1TilgbVDjGU6CoAJQeeEOMfGX1ZmiwkSi4YvK4OVLU5v
TSvzIjU3J2x3DZUkudNuzkcH3Tfq8iHjGfJy88cNZOGAU/KQDO/2n8cKup5/uBK2WWQ8VOaSmE0n
u2VMLzKwF0CZgnazdTlVIqzNvMLTLgxBSwxM4ukdO4PMi86bu+PkS6fAqVp2P3/OE+uaDqnqARiD
0ijqvdgXUbz33rpC1AIfH2WL4EkC+iRitEjRPrXnEhTlCymqGND23dgQtmDsr68E4Tzu645I93VK
O1/Fya9P4A1Z5+GqBrYY79gWQkF8GmhHgUrRA8UrMB3iBsoGhoml1lM3s/01MOMNVhzBtL/CijQ/
3BaawR5bxcDTkuewO2LSZvsb5YF8YBcd/mUHVe0SdU1XteDHo1HitpbwIVM24OQGHjFEiGzAzC7+
bqT/FsFInKpwX9CtLeL1qRPOrJBJSswBlCsAqEfRpeNa4ehGcqmDzG2HEdRwaiHwUeB65qgXcE4T
zycpiInUSgPYSVGtej9tCLG2/LFnNIHIUBKFaNZPtjCgdtUgeMaXEsnCbvKsOin4ury8TWwwoGf2
/dQciUW1N2dK8y3xpUYnvgsW53V3/++PMdX4mVq/MnwOeKvcZNL5gNHpj3By/Y9mADeXY8vPnCJq
JR4FGWm8FsDTqPzg6FVUfW+HJb2HHbmBx/325SEUboeCpbqNROT4GE1an+2Go5qiHPt2ExOxDwKv
l2IwoP0BD0zJgVuQd5GUz3D2DFE8vzVx/H3R3J//cpOvQAbxo3wvu5Agwqtp/qkuvF1n0ilj+2kO
ZZaGHI3/ei6j+F0zTHxkkxpKRDOgXb277XtEQZ5cgVjUYz28BKL3YR7cAxZ7Eqs3N669wSIN7EWd
lC882OH9SRKrr867x+iycG8uOZAT6DVviitwb/uuxFd8ADHmofw93IBdue9vN3ul2xrd7tc/QLB8
TuDfvF0jk+gIl2VQoBapWL5g3YIHHO8s8F45bTBIH1lIzLE2zCZPfR4IiD2rfRR8h9Iy/HC65ivz
mQq+cyaivjYTYxwAesxjPEn9yxFTePklO/QhwXT+qW0aH3hjndx70nxCUJb8v3jeSCv7DMoHabhi
3ZjSXBTgoBsJq9vuEaIfbaTGRHG0n3Fcx7MH88Hwz1ASFt0kMKM7IZggo/N1eSoOGmbuJi53M8cE
srPeeGwOVd9PXRBgHqZ459PgQFmBVR0o1EFcP1ncrbOGguBtWNg5eTGqGp6baV69s7WwmKa9c5Ih
uAKT8ovFSJRqL5f7dlLBIbq3Hw4WUgLj9kfSfmTYpXCovfbAIqZFJTH+rhvzvaN5ElueEdTyVzKW
cl4cmMiLHT3EimRZ2OR8/IDmYIAswh+qEnssiXoemekJkS6k4y4/vUzq/NRWpqyjPqCKq9/isVcm
oBD4KG1mIG6noEKbWrAm/avZ5bb90g2GmVdgpDDCd8hZsN7qUlRRBOJ/tgslXwum3Xo25JKNPq6S
NQHSFSLxzGufMCmljvJI4ghsYfObqpZ0af+KTAKm8sImf4PLNPgnqQXcGniWxIfPrcxYm8QGkscB
cB5p1rO+SqbYgVwhyIbTm/wCoP06L1TWJf/g8x2FpFxpwVdrnClD3iUeCG7NoR8BED2n2Bl5C15D
knRodpyYjdRSjvcYxTWRItFBiqwou6VolVPjymfqA6xhRtzPIB9gvuZa0ySoKCWbjYnI8QiZCZW8
BJSDr55FSVt7db2VlK1beIhxehJAuiD9ANLrxuef+0KFiF1eoOIp1dOeiNrGfqC0UVLZ03ofRbFd
ygCafHF75WchLWYv14CWwELFYWO/pTe7gFMVJv/uQuI3UiGsSiQ63lDP95ldlGnbzGfac0RhnCIW
wSLmttC5VQtHiJ96SnDjDJoBx5yWkDA1AfGdqCF0CSpzl5hN60PVqbRCDyNYOY3Vb0GLDzAWJW4y
1TRFZB4ssRtM3D13Dt+z7wg+sd24wFbOqPUep9kIUbzkEsBdKhX56sojPURYBmsxt+fUCl1FvetL
/slR1rNbzYank78aviik0NUeTFCHozY7o1AHZ6YqE3nLhArdAbTqrEwEHVsc/yKuuArhoO9dPlBz
49w9I865Y1Sjertjh+Lz5th7t4ZXWq8pKgWOQX+TxZa3ykjPKTrUlYADbq35e2f5sL8dChdMf99f
cz6p3L9e+oKb1U6+m1WZYXwb5b3qk/KCFRPEDiuNRcg8XnTBPequ9436poAWIoLaJcM/rI5GACvm
n6uU1xTdrmsXZyXhssotoTWvfCs+7rzc8LpUCUVACB1TAg1LOso/n3qAGVFjVSx7IZL1QJfHg5zV
qVdpvqUCTh6wlMxTKUCimBsmmDSswRF4rDFbquTRpi0T/+E5rxhhF4HNZIhgaA3ZEAnUxPPGkJOB
baUYN6ei2YL7K2F+jx8tWSzvvCnpCYU89Nkx4J7lLRtyvjdXIqU0fwf6EcRtMWHq3JqhTaYkNVQM
PaDEgDf5+dgaTYJNRnrPyBIn4v+F/56Z0K7ZBwm6uHSXvQiHorl+2jnglDhW/AX5BwW/JP6X7sNK
+w5Suy0DEUu8WDiBL1aJbzqVxqkGZuQL5j++dz51hZbZ8zIWKMDSYeeCN5k+3Bz22Y7qy89QJpOz
LanDxXMjhvGtxlvTsnKkWb0LMOasSQWgYai481Lpf1uaBHF4XtqvrI9As/JAGE67tyIFfyLRggXL
b7R5KxYHsneWx7FUoZUcnq0kZZczDau9qh0cD7HHpsIygOnZz4IrMHt6cv13H44/LRusgua9fXZu
vYn94tmB7MsP2WXq4yxgXgDBmx4WzB0h5ZP/BUd+VE5v2LXx7r9+Eo5pmf9lQ90yhSjpN6q5xYra
u7kJjLwPuJ7R+iFJ7S+rq9V2OGiHJJUDtJ/u/vKIHpu9Pw7exXUEZ016E+Sx94RDR+l05fZmXZBW
DHvIutS9nOdatKQ2n/ytdI2LXI/t/ZTfNrmbHe0pz37zPeb6w2oFf0JNXC1u5jrIYaNZNNNFOzpS
MaIyVY1i8cIQXFX/U11zIs00XObzVnWQCaajd3D7bWU6NFnj6SI8+Wr9uivrGv/Z6a1eXvp2NN8F
9NlGlSt8bjy1UjIuezKoSXh1kGdZirrQgsyqDCqRiH9OZljPRlUdqpi0ccUYdvCzzjQrqrTk02w7
yJ2Oy3QREFrww4KPTfNFTGuk3SbZCdjIMTPO/aWtl9afrnRDlCR7FrQZdlg+DEKL9sVarzQcLOBa
LTdiP2n9BjzSuaWq6RXwtALYrnWvjQJYEk+X2C9aXDuAcr3ycIo7J5F9vPsjzZfYIR04pV2WNu0H
auya3mPZzKzlt0M3jXMXW+S/4pibF99kEvpPGGyqUWPrpKGNZhpDKDq4Es6efW2FhjcUrsipfXw4
eqzeDJATc1K4O7xiq0NwtMOgYEGTc27tmbDq9EAwTGpI5T2iy7mf5UgfUgy5InbAmg9NNmkYXuDg
BT0tw2PIa9G77Nlre3OFuI+CrPS4UeMFLQY3j80wZlmJlSh9lfIBgon0aoLHWu010yo+44UAZ7E0
6PGsf8JSivwIjcVym0ZJBq8/SLYnhH9RgcoWfA2JNGnAcGLW51BBBsBCduJQOgEG5vHU0z6NnqSm
CtzR0eqOxZsllutqtFUvlFbB82Tzd61013RfC25G0ydHq1fEFkqd8FNd+IF891fQKkmdcbgdWC8W
CE6UMX29q+duzN+AyCtY6ZNjCostUb2m3uZv7d54Rw4IFGvY+zgmz260h6dHgqwUCvK77YYjIx3b
GS0DyDBduVYzeOdjYABvHGGrVB1IBpKmqvOHmXvVSDpYHLBtOR4di7aqR1iva6/VShU1xBAlJl8E
3dYQHVYSj1oeKzOfPgUTOKnD6MRwYiv9jRyYJOkS50QWSbMBiHKUVnQiiBEZEeenNNAngri5uVbE
KUtICQoBOBu5y9vMrN2jHdiV7N6AB6bgS2BDhbxz/UfHyZxqGi5NMbfkzuS7VJg0PzDgyYPWBo+z
C6S5XDw0Uq+WBoC0YVhc07zx9C84CGTukf6/QgBolYSpfzq35dOwTJrC+io7l8PIY9M67RvkXpyg
j2KFY//DcmfpxkMuatighZxrFZoEZL9VWlb7r+CxQKW7zBerj3T3f48MH/0HvTulS/nq7ZgapA8V
8IiffjSnAdQaIMvEStlwqudc/Bl8bw61cr36N49dih7AGpo5RCROW8yef+yhCVNhMEs26rzvc8dc
TOVlxH75Z+zB+jDfMp+ifRrr29bekFnr0boX2dAWvmgmp7X15Nbu8suio6zt5irAkKRmDXibD4AT
isrxX7sbk/HuZRbQ0ladSjz7y2XpD9l7gHB28ci68BnC7L9YDTbP23mrfoA/N6oF5mft1smdTzCl
GM8Hhc7tnB0Nx8mrIXjoPPHw1X0qWhUt0j/4llQdGAhxg0jGgPV0+W4HcCGyt6LsLzzUp10Qk8TL
bHY1JFLaQ2ofRHKYzTj7TONXVCPk91qxULmca5STtFn8szB1GN4WR6YYL365QQTQglNnbPHE+Mvw
NVm2LtV2aNA/SOhDXkqN+F9k4PD7EY8pSE4l/IO4OmhAsN2EYhPCyuuZvDdy1AP2IMvpN8oG7EKO
SkqT4FTV9gNmBABRt/ZNUfJAH4fgdG0BtBxqEP8Ygsggna+dP5HyJScHMgg9lU3aFFkk4Tb/Jpm6
+iXEgkRjnm1C0X7HoJhXPXYbt9EueoipDW7OcqmFjWkWj20qGCjQ/iGXIDUrDpbjO6iFL26G84BZ
t7RsycqcBsodLzQh3/jNCd35QbwsyLsiJi81IlTos1FZTkk9JD6KQc5gcE4SUh5/lVk/VM+OxyqS
8s7Sjz4XImLPgTGVU7vjXS1cUv08hniSndZXulkj4/JlfYgjuH4Af293HbPcuQLKrxqxJawSR4TI
IMnvjTwtpiH5yf5Vt2glU7uz8uCWSbReW3Hcx1uf3slx98MtFM/zsx2fXQUA+4Gime1G88Ake6sS
CCpvhW6cNhiSiRr/IY+M1zjGlXpI37s1VSFUat7+l7+L3LH7r1cb1r73CwDy+6mJfJFX+J0/VNfo
yW7rDGcOelx5cO73dtXAnDHUCoT2SU1FGHzSpbzlLx7muG4FSUNY/fv13RopFmZjqhXAtFSb9Pfv
rH2rl0u26K7MZV3d5uGiGZmdAHhoXAISfp839uMKv1fejOCO9+DjwdDcGHkD2xpXZH0voRTLKpsW
L/R72XU3QbXKRUKCr11o3PmjK36LXABawuhnZy56Cb+1LlyU4/qpAeaYGGOH22W/soE3pPoGfvD4
qvZrsXlziR3qJJSJFYEGZABPtOXx6tigi6cW/YBkmoj+U3gDDwfYGlQ+tDG2u7rdvxdqVoT2eq9h
Lj/mVh+A3/4y8+Kr3RJsBAzR3akunkT0+YeMEvU9D2npOErZiQuz/qcHTuTwzHW8FNYSuhHfiC4k
/LPy4wwVpcGbvgGpwtDB6pm1aPyGw5NY5W712TigcADZBCLV5aI0pAdoPWvBCVqUxJjicEsxCZl1
WSM2kFU6oLbP/0+E6mqbKr1hpSmzHEyqBKN73ayVk+Ufk44TDj28jT1qYgL3Uc8vmBBynDGrj7dk
O4pjfgFmbw5dFBd3ZarBSlM4k5WjO+wWR3BXKo+elxLiekJD7lDJB8mjeh2a5NG4vSdtovs+9WyA
TAdBYb8L32fiidNa6agNQHOpS67pRFOnakuNBnmBg1uxDjeZjQgbKTeF/KDX163BQ/IKf6xBg+5K
DuWmtYRUZBlljCiNXvQKZ+KJpk2CKsWesTxalWwoWOmQdL3avzfP8ElCftPH6j5OwQ6Gpo9muEFG
Udx2g8jh8b7I3SiFySXexFbG2+zUMg6/6udtn9BRCeuTtZCXi9Zjjfw1/Zvpv65bU1fFYaAiSWh9
pIprSjaeh2NLvCLYoHv9HhUBywXyQ4EpOxjPEBKet9O+yfoRsbxzXUg7v8dFGjf7ACFYv4FhRRTP
aOi0omtDeuf6ZMoaUFitvn9+rUJSw96jUEoLsLeD+zWNUczrIoW9lioniB5QVPmSCvjizD+ggOP/
u0XxvwyALt4UwVZok5U0bdS1OUsw2gdRPcan4cehVPebmGk4S/jVWyYXCMV+GIqyT6FFpUcRvfRx
nGkSfzPQ/dkAJ55hJ77khlGklY80uXxG5yFqdtApnPEzCtf8YXjFrJDeWzOwEwYIL0khQ+P1DsS/
ndu63MY+eftSN+prguX2IGpFROMU0KXE9u79m9Y3TKovEhkmQ4K8GvgXoKcYVVVG546IJ4cTRWbH
n/ApuszjOVmYdvpQ0cNjMQ3iVS9CJjm2R0Ewej9CgrdrJmjWu8yOYm3noaJVMNmLrYGCa3mcvndi
oqHv+EFjLYiGRyomH9Q9hg5t3xBWRf4rEPoRpFXGoFxOUeTb+G0NYsI7eRzgMjoCAwisKYN6jOZf
jcwK5mj66vdktgxgJcJTW/2+cCQtO6odngSNcvOev3umbsYLpFw0C+GEor/1xI/UKkVP3zYZuVzU
qSM1Gqz8HkUj0Dx5HeOvtOrJbV3A0KiXAEKjuW0KW+myI1bv9yHKPJ8bVd6rwyf+StJ+K2w4b73e
/wFyHRcBTBYHhf2u2kEOXXYkzooeCrDLtsV+ehTWOY/hDDsVI1sFm6fFtrtqQOmXZtBYDiBS0EsV
HZcMoc7rzjoTx860VZQj+fPJF6nZsFDi9WNy41UGZCDypgp1lFBbGCZFntjU5vuSWeNAersb/kwj
Q7uwQ68fgpLd78zBE1nAF0uH8NiGSWh75ByLtxOqmEulcXTQhRtqCVc2G3WHnW89ICk3lV3DqiAO
b+5Ry4NG0s0tiMbvIZlGd1aAngQAqmYtd908LqCqlI6AYA0Qkh92U+HJ0ZxaKF04OMLjV9wqVJgM
b7nJA0NuVGsO6GTI16cmsm8+eanLbtrPzOVQfYtXLHQ2saBiDn17SjH2QuB7ARizs7oJ6NLYoqXo
wsOAHVCOBwzfPUMnmAXH+oRvZ6t20oDya5FcK/J1ozF8+P1V/UP0+AuYGcGPZuckVevYYUURunLo
S/ylylC/awEINkIv49tr3m7KTHSccrziFCGmlVS9+BqtFYy6+LaLC/AReXLH79C03t07u6nEw/fy
Zf4XM3r3FjAKGyVE0XVs9ki0St3QJ/fPklCrlhnuwD1N0jC82asJAz3xxK3MxZ1D9c+geznKjodI
SapzuCSjfpKxrDj8xeUeiYTRgj8YexyBF0Lhi/SenWLE/aElQBRh4Zp2Oh4MMOboxOKuBDwpHnYg
rgzrBm+teFSkcwDE49fxWN41MXnKiJqbJ7ZmgERN6t5PDxcps450MliVhWp/0wAk91STnRs1X2Zn
MAdoZBkNANoXSPXUCdeUXaeqPUdvw1Wm5OCXevB5pEXrpuvezGh3EQ/RRoUCp9t5mmzevJmCSV6+
DuzPcQq/slzlVtyZd6Prv7nZfN7zLPZYbESgPWHr2DYbTL3nWJ4tJ56CQJ3u/RnDDWQNuTdhJ7Jz
TDtd3Bsx8tr3pT3ZYhn7QCEz6atk7S405CHUzcl6IDZ5g/y9lXcy3g+N5ACHImiJob4tmI8SXtpI
xSXR8wsSRsTb0jIDouZ7ux+TnxvIT/3YRXXhI+O50vc8vRBWW6WzwXPU8RiT/bnnayEP15ursOpS
LpIOqKXh0Mfnq7tRwOXJLnPw0NGqekyFYVmoz9XfSvKSYws/iXovcLt3RjYyTmFw17Q07PnV3rJw
/GgTtNRDigwb3TwdLkrIaUPVJIUAi5qufhvmXZ3s9dcUM7qPEC2RONt3Z29/Z3fgC5re53k0FTNe
Yll7f0vUIF3D76ym2SD3DiBzUcaskO7KuPWz8gXQV/jUDUifdhMcdFIEZKMsgpuCj0H1X3JJUNOQ
Hu9crGBUlvQwViI0oYvj32pz0WlHXpIOn0XC6rU5k0QrWJfVaCSkO65fLacjR4y8TpelaNhdQSzo
8I9WbkAA/tcGjYFa4Ip9iir0upNV2rIVUec1npRdnhqzzop3YZ67C1oI0tNzx82h42Iq5CUNDDX2
MNpDX4dcWdpt+O+mUgVMijjnct/KPVAqp/4bY7fCekk1Zrq9R4ZHntfQOxSfhM13jPrAD69UkQ9s
TBWx7r4LXlbsTOxa68EIiRq5o0jYajCRCl+3s7ZlWCLBvoZ1w6IVvxGzAxd33tp2UFRErvrsclhR
1QJsKF5k9EvO6WQ68LSA4Q+dHL1Eiys83jubC+LFld8+Bi1FzrdxIeveNX93w/f/KFmZ8MkEaVo7
SXqlrbOMkIgiPFr0Z4OGE+W/Wsz6niKLjraibicw5CTm3SQKdjSlsiaiADy8omvp0jEifYO9bZYE
I2aAoBrxTT6sDjp/FY7YTAlgWGI3s1Y28o33qEIGDkSZqHaSa4NgMT2lItjoHeMbmBWb5wBeunj7
LLa8HZShysvopbZPpoIT8YQSZaH8Ae2ZTNxbDGIIyk+L7Rq7so7bF2xUDnCXt/V2TUhh5F1gh6g2
QcXyIuoLFTLbKI7kIX39M/J4J10RcimNc664pyS0k8azevyr3RzyrMDKtNgrEWNZ5B8p0aYQV6vX
Pfqt8oEuKrmT4YZVxwpvpJY9JrE+U69+Q5GMPuj4A28upV2BtTTw/FvU5IA5vpIhG5RExRFukGOm
iuHYtw1ZBo3TDzC8EMU2GQjhPVcgYXz9Y7xXFUSny6wY5PqsZv+PgrxaJs/X85EdEfwhPBTgOOeP
be0ZXeG0kIQ7GO6SXTRyuASCX/yKyjJy+7u9IkJEKjJD3sOV1yTH22lYcO7ltfUvw1v1T0j7Xli5
goqQ8Znjme5NRVd11g7r+7qhzJF+XZwq5NFBAufGiZx9b/+tBBKj9lxegFwff/ctEV3MydKFblme
ObWKCq8sr+Ripz9lucBPzOa8U7z4ZjdzP/rso7TVhYLPrTBh4kG1WhL19+k67R66dtnaji+uHkEt
nIOaoJz3LfdvKPRO/5/HnqNLU2cxjv9ujOmVZMVqOP1l4sx//gHxuy9MdnNQjUfaKW5yvms7Ds2w
bH8bET0z3sZfgZmSdlJltr56tJ9DbiZpge5RWDhOLgP2gvkPVU2wQrg49fCG3gSedXWHVx29cBgx
WRm7G1OnF13GebhJvrKVVyO1tEkAhQuCKd5zc3USieDYkfpWTpKhQYKF8km6heQVWglmax/lob0T
e9EL6Z0aKnbFiPo62eKGoZudy67ANpJca39Nvj9mjF6HKufQeWQmQiA33rMNXh/jc28s5R8k2F4K
vICIwOux0aBOnFpCPc+C20+aUQHHnLV3a/bwSj+Z19l9tDEqcvGOCRNFrNyNFcf2aG+3tFBUbgK1
tkQ0THtdHQqUYig8eMnqJUMXaJzP9pAfnevmWwhNlrp1KzsR2ojb2pe40mdqkjdevjVJvSYlGnzL
9dzn092X4nohXsHb0LpaSYGjib+XsPkbxJjcbmwvMAnT8RVfBP5AIONGZdCuffmCgqYzdg2yNqjs
LMzF0MQ3tmlUBxp+pYSddMj0oaalOV62J8hUDYzop7aDwn4TVNGZN2SJEq6HSoLTve/3wyDIQPnx
1iAekCLRyRYzJ1/EHfv6nZrgJg1HRi1Sr0KmhIqvtaZeCREKAzZtxWWZKDZF6Kq2vrMUARC7YUV6
ew8fzvVMOq2hno0r+aZZx0nG+NWC/gjZox7/cs7iPxXQhjcUPhRdaEb+uAN/u7OKhSzq8K5UEX1W
rFSrSu0a9IXUXHkMk8qVHF8TE40a1NZPHr21kW0PisF0paMwVbV7b/muC8NmyU1sGOTSAcGpi0J5
AKBEAoNTE3nLOxtGf+hRLN1zWH3FlHLwR7FxK7Y15k/6FUEEdULyx7l9JctQsINVt2C8iS+Ayp6N
/HopQEGqUuKX7pXdCpaADXlmXA6xk94YWzvwaJnEJ7+oaFQhvK93QgWMlrkWgEiijU7PdZAYJVHb
kddN8K41PyEN5HJcHi9bWKSVB7m3C8YZ2pJcvI7f6DcGIeFY0OPe3jE+CfYRZ0gll33kT2M45rXk
ikU0zMqmOuJVr5+v7bPbsSfklLDThinvDvgWAzr65UYgBEETOTT/GeRkGoL+rYBJccUH3NvukDDQ
Ozaqkmi2Vfs418n15kqFp2i4yhMk9OFoWKCdg1BvYxVagc4PdZiw3bmRzoqxSFoC5v0TIO1SFuRr
GL67n3GbRO0ihGbNMNOI1UDGlQHxfi30nkgCbEVAYyN4zLnRhOGj7a2k2j29dS2bF7FqRA5pTS97
TwJbUENmtJTHGtjAjv8Qi11S7qRT3zBfkIo4vD1dSW0Sp6zhAvzvpuIkdvQYbzkkyjJlH/fn9fhq
9Sr7ZBSP1fGHTHskAGYbc6yQFEv76N3x/nqtgrGXzU8pC4f2phrGcj5PEJBScNuGMPUoqN4xlAZ9
6na/wjIlrNiSyuPNnAkQZNpRirbk6ej1zOv6bO3mm4Q1I3Wsnky+JdTtU6lBUiZDs7ZLPdIfzJ3s
HLA9v3+8BqZ5f/oGpUHdQ5XoCpAmZHQnumgm8P4YPyo88D1XLCfJPfXCzIF4UQJ1+MCREdXQUXma
HKni66RuP1SPJdLAOErT3WAOdNq0DsWlrUsxYCiBkVlr4ISiicCMuI/LkCtpaYG+pWdfj3/xFKx2
g2GrMwR+JD4K4ER6Og5TqQzwyi7uHWn7tMKXnj9lj1xTzBRLJxJSYRV3Ea/n1CRw/oke/p7PgMeb
zc/AnRZzNvmDflKSYt70C/uxaB7NlTAL86v6DvetFNGDc14CqxAdMCgQuSIq8/flUIKn+TW5Uox9
AYgYpLX455DR/0kuTgRk9HW9ESjQGslpkRhVKAIy3saXNk2tEqH2aXVdhDO+gPQbkTdD/xnGNoEd
xy97kfu6Ci5Xad4pdbFCsJIvDppEuSVMcLQsBXWNdOUvkX9kPKkhEb/ZEvuN3Mm7Dxfr4hPZSwuj
rSkNuu4ZsLjt/S9VoL7bTCjgcdJMbLtSMZvh3dxQm6cHsEOp17ur69T/ymwdMSwnq1WyZXehxW4V
8X6CYEJPJFYTl58Wb3z863ZGodSNgggcD+iiwpib46bMoRLQO6yoQpDv/Ib9XKS2Zz3X6RYfQuQs
dS2uDwwi+yWqz4FFTj6pYmbklcL6XmFe8ZwlPwDWZvQel8wPzu+jiiW82xyk4G5Fmg5fD+kv5XXf
Wk/ZhHpCD1K66d6eAMHw8OxSZo32U13D+ccWxZ6QulnNxlWovrnk3LZB2nLspzXbB7mPXG5ASk0C
Sdmb2bK0+N24vDLF2qyOCCwubHwabNQAPBUdtsKiEwbsSMEwraFFm0qQD0sRH4m4px2hKpf7UKY1
/krP93a4aGWWWYqUk/S6N50hNfV3adtQI4NQD48MS210jULR9vtqfxpgBRWYLxtULmr6VaD+r9uz
Ex8vkL85mXoeCZbc9Rq7yCxxYBjittOuyl1P8ze8e4sQi9gwN6ZPIHOu16Bk/Vukwke9oHZFbag5
Di/VQkbr/pULmLCOBAYh/ezVMUIzT4EDVweIt2CposgeL+kw/w8uDIvRjqEWgdG4jpT9Vx0kwoS6
VILsdZ7ZwlvyHAEt9CdtU+I/upFuCqW3C3EmvGGwfT5cXbDkJl/uSdnaxNAgl3qcnhnqjTP0yhU1
DOt+eg8njwgcuO2QNmUO1XL2wmT3ujsohNmTZA9por6YmezXvgyX39WniZkhF9DEQw+Nedcn+7er
i6zxDenO2i5kQbjiuXIUdVDZCafMMI5Aboo8WDzXAy8ul2vRotz993Tl1RBDfe4qdroFbavG4fZS
XSh/I8mHGd7pSShezowtGy4K1sLFf1OdjXoemk0MF2SlUUztX4pzmQmvWUe6cStWlC6C30ygofpI
PNVk6/VKPTrmDByd+sk07r1A1dtAuNs4c19GGsLXhFyCBBOg9sJ/sZzXS8+T51wu5xQb+qUQWWcf
icEO9lvgmHqxceSv7yD8Vn/KPX17bb9lgsuXr0y5lNmwvxW7FllHbugs3Bwrfdnlw//R0QjxXLYg
lNKv0PVGxwfyuHlcuaTgvReeIFEd/UExuFthjacVSzsfInMSEu2ULRydni5c/+e9IdSSQqaBtSkX
qP6ybAHgfRAu82/gPSd/USt2LjZ48sW3DtWr30oREVzQAnOejSuXSLSAAiaSVZdxNrsevSdFZRC1
Rh/ynZbxsM998oax5FmaFxqyqj8czJprlxE5/4WBqZhspeyhcbqIhCS4qi4e5oOYygYvMUEDVq96
LxVJ/pcrnBBpvnH2xTMGWW3tNOum95uiB3kgTmBS33lJzFcVhj3yoNY/DBFjcoLJr1nU+EGroVPL
TO0CuZXoYReLRuXLw5Pg0iSXuLNM3FWulcfZydn1ysddTHotha1ua1kot1bppWMSL9IBb/6ipVwJ
VfyoKIIBXLCEDdEfje1xcsVxpjLk+WwBJUaHaVGiJx61m9c4kc4pt8u11CgcueWd5CLMlJ1kiwUQ
VzKo5YMhOJn0bSfMXqdKtL+XT1bw71g2eAZbyPgrv7pEfifPmKZhfKYXnAr/YE2AfL05ycZnCvEl
JYifzXk44WdtNO+r9pgQizg6sfn8gsa9rqc3kXkHHycgzQtO+17zg4/MYh5Iwe0F7/5J5GSpx1NR
cidRIRC1rr8lww9L7dAMWN7OQeUmbM18HTnwAOwe7jT4UVZZtUXcRwJuTRMuid4n3xU6waOgTCeK
CgZAOP7/6ORMS6qdnwgTCWUlZ+G/zUYDbscpLJUnAqH6pSoBd49Z/NfYeDCetAQPnv7mTurKHvRW
Kiv0mZZTUuAvkXhbkSrSEvQCjXrCUrZPwzx13ZCAabtgGDa/FJbl9g8CSz48XwjzbTA9pfEqCGaf
jz6zbN9U5ID2G6zgxcCGZaZabSmspSU03fl9RV6mKPb5NxTVykQiEMbSmxXxnpYUcgYPA6JvXc4Z
IUgJdJlKndVtIEk5lqTlVwLDzzZ1FL3iY9YEUB4efQsZzNQW1LAg3+QJX2C1rwhcUutg90WUEv8J
KEwxXULz7eJOWl+v0lry9CSBhLhmd0Xb0qfyCSxZ2jl8PuU+Lrx4FljsX+Jq99f2qSPKlnbXO0+g
OOaIAbXkYd//PAAn/LNQ6SJ4fiDfnClYxyNrEjY55YiUpQSwABCwT0GkBVJkQqFaRnUfzLFswE9V
CUwqIgBMZwt+OE0QGE1J4jBwirTX28RQlstfSGcBXXAqQXR1TuRbwicYCfovk/KkDHMUw/tNw1ti
o1A6NNUr1414wUhiOSChx3bO+ec26232NS3toP0KR4KkJLykIfcQ7zNOfDMR7MttW0Vs3OLuW00s
Qiq2fEo7nQFHzWHLVXEDggIcXwE8EsISISromGK7icMCfQ2srAGLA4Z30/MVQMu5serG6HD115fs
9kysUT8bYv2JSmqRuNtV60z3SNQGHAAluF9EgmRxwNIVdeMuoZdzQ7qKwDZM9LMEs0B5kUzf2stV
kqqt9qSGWWH53pB86RrEh+JRoT6UcTe5+meQfDZlSFDPntSkFGUnkQEzxBs4LkivyMTTq6OJMR86
HVxoDWYfSyKPgB4ln1+r0UCtcstq+W7/u/4vqGZt1jd9wxoja2W/UpyC+hpzpJ1i1zt1NQPQ3XmM
zPYpeaqe6jGlEt7k4Y4Yhf3OAZqEvQXqZWc5vloD4E7uga9zad/EQl4GC4Bh1KH/jtx1C7rCLImb
NixbOZFbkFADqrtDOCWzK+HqMjP7hQj/S0I0uB8DOM4vTv1z5C2dgLBsBSdhO+I9V0eYA25tOriH
DbMTNP1sWIBWdMWdDRoZKUDE6ZDbIAWM4siapH1j4M+FpPRg9VJ3YkU+aZEjxHY8tHeB0C9Lb7ZC
FnA6j++/CXk5BGJo096L6j5csKS2R21oDKKcW+HH2MoXhrG3I7bjsqj2fOOjMy2cQUOGyRM6KETL
5wC4Sh/+TU1rqsAM2L5FlJc6EcOKgjMYVcO3ThS1kd7JFvp9wUCSe+7AkFH8l1eKTlP7WYWgmW/G
u7ZAW9FWcYi0Xai4PHygVZTy/87CaYEaY6XAcMYniWNEnZ0flLXBM2JURFQuSHmzk1GtvXBEBJhY
sGPrJ+dykwMu+Jt6ojrSyMjJsM+rushrvLoQLkL9CAQxPtUOzseHs5XRHg2wf619SN7CiGJQhhDk
yDOpu2YZLibva9xtuBlGj+UfwrkJW+hrWZm/pVAodxsPK11Emu3NYv3qHfAKyRcUujCgqHAofeEZ
Vtb3z8baes2Pdx5AUuIaVmIGuAGq5DeRQCh1JxoESyDYycdnWplVV4t+9LLLiRzKC1FrSvTWESdH
WT/62HA+JQuo6eXVorFVG9vtdgdhg+a5z/dW2CzkxR6+VpUfkMz0qyQLoMr+HzKdwzD+4rUGDYvJ
/YMzRHdm7kxWyKfj2hbKrxiFcldKAbzmGPOXnxZnKK4E6PfwZrtHUPITox4HYSQ6IwQ3plEKYLzG
MeFKGIVR9VjCvLejzIz+kpQ0tp2GpnkC3JsbONlILtF515CFvAvaAFo5LE0c/NIE+AAf/+CnqUhI
bnWh3Z862Po1cPLYKjyLGph6H5MQ+wpnb/znGPqlG6gKwoXADIwT9KvBYR1xuNOSuvDIbsgTBVdh
LDDQIFrK4o3/vaq2uKEsI4m9lqzX4qQDqGFBbPI4igyI1i31BkkeODhUx8xFo7eeQhvMTRMoBNIK
O19hVy8ZQHUaltd4znet+JFy4hM6LoKxj7YaGgBYA48YxUmxIGVth/W/iMQtdcyMmWOfw6VBJnUk
5ZN607NF35WaKW39q4TCOIBZDGVzxw7sI8ZAc1KOsGDmanjxFxiAPrL2Z6VfdzJ5TBX0ZzkD+ou5
TOp1uIMJI0v0zlXmjZNah2YcFMRLOLU7MdR14rPiHBWZEALRRycLoK+7E4HiVEXjPA7x/wCJc2vi
5r/oRuBooEcA45akhHQNB7/pBly47oumn/rtjz5R4rs0AyUD7rBmsl3eXqmtJr+YPSRYxJkCaBpy
qTzUSh6jxWv2JheYkd6GLaja9A2plfq/vyt8E9MtcMGgzIsp8Agx16wWKTOtb/ugd/mdnAp80ZK6
iTOeVS4WjH3jI8s5jCUoHof1tjWcq0oadeDnzJm8kdfyX0RE1Q1NQWG3QkeOVE34IXf0lZb5Ly5/
BXWOe0rFTTezn62D1YlbLAQ/Uq9r58j0kc7nSegGSoBWADqtGGfP7UsUdX3+rbF/Y/JGPXFJ0/eB
XRVUspnPHl+BP/t+hylXWMzkWHbGv/ieHiPjVOuC5zZKC+hJMLBMTo4x5MElSR1FXDW3wZqAY4Ws
wvFAXjtzmBcDL9QzyfFuvanoTsVhvZMuwS8rSttEsfOWzLJ2WaJep0zh9c1nGf3qrCgmzJu2mGb+
mMgYQkucynIUehCB9Y6MnGDU+F43HItyiZUxBrX1oiK6rCuesxiQCYJnYTokyS2D239Tpraz6+y1
fDbcNtyM/cD/t74JuNugTCqZ0yTxWLiAAERt32O98QGlWIpBGtky2uZRg4QUC1aWg8kFYtD6Jo0w
4AaiE7Bza6zJEmYVKMSoKzRBcSJ/lb2Jo/N0BlB67MsU8/yJYZf2lTN7w7+/SS1W6/0eXz7NxWFP
RA208gz2P2pl68s1J/AsCFYAEIDK9FHYRkJmufL0caRHiVoeRuVxW8qVqqb//Y5C58kvtkTmeetC
3ldq3FI5EyHKYd40UoiJSn+CKgCDvExqzW4eXkXEk0Dxqlg19G0d2TgFMm+eEkEcOp9FPc9yRMg6
22NjxgjnYtdOFUiM3Bl+gQumjEyHEc2Xcoa+yGhvo1EBrqV5bbHneIE0gu7UrTboNIWWTndNYKpT
LC5a26MLrwnlu8M1u33FoJhkPy4xscgb2Pds9LZEgFuzahyIsxAl9mwmNlI9TCejjy7rNUCITXtk
UbMmb1GWW6260qqX0FNGalZEqbIlmbqQglH6sni3qx2h/7vfM9/nThqGdg/+H7wQPD+sL2/LAtI8
optuKqR/f3ga2f189YzDzoMKLr9PXMaiZmT/JAOXAz4oi6AKKk1AP6HKxe8b+Y0d0MbX4qJjFGpD
ERpQSkHJfK8vqpDPjbD/5/l9d1HHh8o4DyribzkK4GXp+FtAhD3neXVkoeXldKsOqh7YjZWNxC8F
NBdy6IALvqOtwWBnsLfZxlo3YZJOF8dajTMhjORw9dHBpwviJAMj0p9RWg/U/qkYBlyBDBhuWk5M
06Qe5O16kmC71QvQx6iCQIpuCIwQJSPMIqKbavb/r9PcNRl3XU8Wuq66Kot9fblPUHzil8+DaZ6n
JSx610+7H42kxjMtJFTJiSP8RJqj8ZRnJn0N0/uRnm41NJ3oCoL15298BKCaDWnatR0XeFQomEjC
eeDuVudjJql2xEWkCuE2qIgixrB7igSP16Ivv7b51vv+2CnHRAqlbWJfon+EjzhzrYqOWdauApot
fUqmBvs5p6PlXP0xxWaRH2EVsLFg3f3psLLcJBqiuDas4d5O3gVlbM9fBLTjKaOXHfSRp5OXc+rW
trcUSNSQEZUHAuMDoOK8wPWqhcn914lM6hG/cBwzKlcbCTshkC6U7xvcmmK0ztsVcZkRNIp0hagr
U/r7C/DFNuOlx3fCOY4YUXYgW6Nkaq0qz+azrl1ElxFC3oy0HA4YbDNb+RPuVI4ndc7z4uvYAOoB
skf6mdxFRz1Surhq2ReVZ23fGM+9oeaZRXwIG8c0nGeYfyJ8C1av7p/rYTWbELR+YbV11FOry4nV
CaOTWaeliJtwp91EH3PeG8UXNvBmI3fw7arreRG0elxGz1CHmKEuhIL36ixQQEBG+n7pmRXlDVXE
wtKS5jroVXITMR6qiP5tvKf9LjVqZaNxzfI7IwRjAyLgTYMp4nXl7oFcz9UYmUljkKdh5BDvGh7p
Bs+VJRtF3Bj/C+jngyG61ron6mcMQVvBOJ/Lz2maodrRHcmZiN7we+AY9UgE8QNDswAs1MoQVFYj
bg/IRJYJr4Hr9+v67ZY/TyWfHxiISZMX/DzkQb0pNbvoqK0ZcASWSviDtKJaZa4auLq9uOxARyXj
r+Nj8H6/PHPls7QxetHljDLOJT6zrw20YVn7m7HFdfOhgyAqcWK197BApkrLxyT46+NepxLvBUGP
wwwsAZkLwZjNQC1WaEH3igohIClx2sgyNx48NoRrz28YvhBmuXrZ9eg84H8yVOrI3U2wghR9SHVq
DzreXe4ZfuXk22uRWQzOTiKOpJ/ek/FWWrA+HkwNGIWVArMyNc16ri7bBdYyySJWy8dZx/m/y2Ru
vW4FQoR9w9tfN5UizooaY8FJitSHPi7+icvOclu/YPJHdBc8nAim/vUg6ozihd0wZu6RiNPQOgI9
ULIx2OW2q0v1wpmtniT05tIS4lFeJ6DS8fR0N1TGbUO0HSCMswLwhR7oWnBq47CYVGO3hIQ43ZMt
9ORPAXjAynw4AEcrMGIRkyJqa7YpL50MRu/SbAsxkls7sVShOCl26Sq78x8hiagsPNi47alUH12K
gqBwL7OfHfa8GTTdEEq6P/N/XX0MtqOLG83cwHZl1GADRHBDfnBEOVjLCzpqxjICPf0xQTyvvIZw
j5A9V1936cEL6SNRnJWw8XZZ91mu01M8YAV8ESfvhy3nRvNe4cM/xYmpWRgh34dPd18hP4X5JsH9
N8riwcJpbNWnuRljw1zGeKeJR3iXKUAjHCHHhM/sPJZZx7mGq8WuVeTCAWZoNYK7Cv1zfi8+Qt+h
VIdBSSWPgws3plN6RP1lmXVHcr6wHgV/Y2tjF0Gd2NO+B0K6uesMqg6qGgoxdUOFngmyP5H/QL/z
LV+22PwGAveYykkocce8K8oBzuojDyuFuflOHBTrLyp1+iNoBm74qnWKn7RHMzRLCEGAhNCdshO0
fDVTC3HiBDDKHPi2LHQRqiBtuAQRYxDRh/hDfYxPu5s4pfkmw5OIKwPhxrP5tpnnND+dZqyoHzZE
I1adBzpD5Gk/g25mwBXz+Qdr7RSNMCuD+Os4PypiEvnqxSzGxkMJ8lKPdqdbxR6uGh/b/0G+heTp
p2XXajTbqMAI9YhiK3nEvKeu0gekbQDoQedJ4jJYe6DnoQBbVLVp1oPDuktOIhCcaIjuLnoS8JLM
SiZnqU2HQMQbl0uJ6YX5e8Bc7yhEL6pTdlcRwSQKOct15ofst0Q2VshyZdYB4ii+hmcpf1KLYE7y
n81HDyaiZuPPzyHEKSXAAVlkJh1AMLtihz6P71GVLZ4iK4z/qfjlsa7vi74Qj1gylgaQSConB1jV
x/zEY5dZRmCIi/vMfpT8PSZ06Qmvv396vRDVMiRa2q5cu9J99tflOgrhtfXy18cJDY9U79MO091N
m/JIxngFKXLWQWBTNKyhLyVR3pGUP0ix12r8Saq+rEBPXdcyEyR71Rn57uHGkgyfW6Qyul/Y0zWX
y9dhCOEGWsWvmj7Y7LVhLMp1N9u3qHJTu27Wt3cGpIDITPKILr6dFsZ1G17+9BnoOciIDdwdT0U3
u+L1aBixLEFkeh7S6i2TKgpGu5+OwHPvIO0tZ+vb+oTTvASjPo4UHFqmVnWp8pL4VfBC+7l/OPDq
hmM1KDzpDleQmhHtLx/o2gJJb9zBSJzHTCXw+gqRuQ4f+Lkowp/cCE+AUd3WJKqulm3U6/I941f9
uWgwFyE79X7f2el7NRHh0oHaSKJW+IWebLONlepsyZVsgFm81NfBVL2AoQLqSEMLjpWyvYVG9cve
2CFsuNb3zLN+6tK6gTeIIrU0mZWb/zdZLQ3cWQvtPG9Uyi0wdkrxKpsy9vPPAXeK7Dw537Y/W5MX
3ir4+XffL7z8B7M98klqu8ATtyVQ+/JHqaU12UJdRyF1G7b7eWOa9e+5AdXtQrA0k9Am8KYyiZdp
CCEXs++TWPF/Uk3Zi3iy8G2ptnJppV33OEtQdMAA/sZitZBy3MbFcUeseEKGxqhL+9UNrlIuRCTX
e7VlyOKo9MrHWyLbAa9bvvEGOpEgogf1h+lhPN+0H3T4yRbWDBHlBOeUIFqUqNP8ammYNuCH1dmp
2e2PtGGuPqidx9rc9fo0EWB/SI7NijRz4a4wjDCk7Q1HWzxiH2ccSeBOw09vxjctHiF5RRPzPQCe
1T2jld/YGUa2s0GiyDwCKe+LzNizaoVmJeIx7vLFWPIOch2GxqkK9KWQSNXifEO4/R5gWMK56kwh
6WICml7ROub7jzKYEg/eII68kUi6w4VMN33GNixm4Cyxu+ZPDk7bvN0mhYkUvx/jvg5H/C4J5nR9
ydiFhXLEyNQrrgc4bpOCuDBoakd+6dhg8vagliF2pp2g+kwrX1E43hOUXepWFCvBCv7HGDHkbisU
5VwmeB/TQpVC521SsVjmezli2958cIyYLOMhd9IZQYCBkH0cc+7PJyvRwGldVR5/qecptYyf7YcP
5r0xUt5pMkoOaYHmSpxY/+8OZWLVOD5PsP5k3gaSC/rK0uQR/eEBC9kgTMSSPisBok/1UFVGHlk+
psOY2VYnnpCO5DbQ06Vl7lCcpeTLr9r5GlO6lXRQswYGJ2BjKsBPXgS4S2id78go1QjBykZl+a7e
8hrdCNWbqdFm3oOY2ppUzwdeoeHP7p8JT4o2it3gO1q5JPw0xBcLVkBJxKBwwkzteDLFiM8HJOfy
N+7cDYOe5kDDrKG6L7fKjb6wZvldnuXLGsSLm4KBUtbHG1Ar8OPUfu+ioOxUu7pMdT7BBFTCRZ22
dHQmxtjLqKpb7Ci9/qCfHTu9ujQSth8fZI/cBVMDa8MK352tuisnDiJYQISQwgB8INPlxOmrsHp3
tM4SopuCsn/Z0VIVxv2/OzAhGl8A1f9i5gmXd3Pe4grGb8pNLZwbpQtrDpPi/O9NpqAbFD3q0GVa
aeEGq+CjgM0nzNYp09B6+6QGRbgw/JHLoZzyFJSRKbQsdRsWf67d1hgIc9PQf7sDnOc15n1Xx7py
fpI6l/rqBg/EaL3iMWb0hs1GJ6EroT867nHqqTIrmko7GYVZ9P6fZuAuhfOOKRtlCWVnac3RH4r9
mEItZKpvhF5/wGxiqid9rQTvIl9u+3c1tZIhB1zZ9FyIa2lpYkH3LZwleohT24/SwP/G37yJHtwM
1mKL6SjOzqkFY6fk9gUfqd5jO6Tn4S2Th6Dxp7IYMJ1p5fTyOONxyGmLFGiE/8BIoNDbRF7RSp0c
duR9sYV409lxIdkPbDJyruqURpXrUqi+Lxl+6E8syIZJN7NUUdxN02tf9l2SYMTZjJ6I8umRT+ua
QVCvNyrmWMNId80Sh2rIo3osjjfkOF96kgAf73nRiE9jXAwBGu21GaQQaqYqoGs6liSDiyr4OB4I
9BwyXp51ZNOmbF0ibjnDIpo8HmKl0uJG7Dr3fF6zH4hpwTXPNdI0KZLj7AgP8U6/0+hTbSWMjkrD
e0WqkZ4iyKdkE3q+6SpnvLXWSp7HW6nxENxJHg49xodc2lN4oXCUhn77K/egYoybTmxJRz9op9Vh
c2dzCXJnreumJE79xeT6+LiXg4sccDhSwYATmpe7hKspAR8vVI01cpPX96pjFT32ekP0/kRSJiqr
u0DpjxGqEJBGykYxjXtYcjnNfWb2JPM71N5cXeaEB8+f2AdtDBj9Fy3e3sYjub/N8YJQAKu6NuAg
GF1xc4rc9r86RAbOlGpu67P+4bOJM9jyrB4pBJ6MUlYTrzsGbWKjb1GtGcOlng1/+QSJJcmaSYze
/oRW6Z91fWsDMw6vhrYY8sw05K2NM/re6oLjELIZL/UmPl3Ksufta2LWuZ9kOhlFm38TcjYJpi1b
3rijXwDRENqClYFwBIxL0hVvWMqf2kXzy5VPYfdt8hLUhNmvOdhyJhBkCXmVySS22V5mLowFDdoH
rNMR6GOnEoUkiVgDkOy+8OIo355uTCaCgB/6Kx6O18rKjZy/suJvgZ9Gblw66XSNSc/MF9d8Pgjr
sdtLh6uZglCG7+MhKb+oUFl9qGkthN8lTyHva3qUOyv3IswRapwLVCxPhaRrAIZ7Gh5ueNS9yKZW
B5GTLtd7O7pGXB4GZ4Fdyx74xUpsY1g2xw2d8Mqy4otCwKpAcVWjBNDnhK2WAFEZQFHSO9g1cMxY
ftDGDrKhsuPHGJWtV7lT8hqRMo9z2+bp2/3HSyrLCIP3bxdaVCMXqLDQCC78a3rbAS5O/7+Rauw7
wIJo6eq07UNHp2ndPK+uY4aktAZutvaOFhhuRd2IK0mT4fl+1uCVfltnhOLBTd+tM8dFvCe+zWm5
uNlbXv9h3FUoCejEJPLSx35j8FZSAZc1ZmNhZDcf3FL9vYlm0W8FN4/OPVaUc7d7dNzCLUjsP1TW
FXXwy89m/j1WDVgnMtJDAjzkEmwJEN/Nx6ajuldS8SEnDKLLqZuZKDjDU1xo7LsmI1k+qFqCt38u
r6ibrGNbpDCEGCQOUpIyhO0VCh+k6dDbM/X/U3BF6+RO1qxd+BFSKssKK3RSGWWuQbi5ORkTHU7n
Fxng8glF41OleXyxPASzcR84IS570Ow97EA4JxFYPG4/9hLUxaNHWSyFZM/gmL/Ozd2MDkp5F+Nv
AXqGWEDsSKaet8yrXqP/ABPIbfJ+FXLKC4lMDH/cCct8g/39bRESZnQ6fiyXpis2Y5c6nkJX+0Je
jA1EilHpLamKwguqtCqfO1Y0RDM2XYvqO5uhCWGmqlJDSh+69YBrHmi7F/6QX9DTof2ofgPOIGWY
aokb6mqRY+fulu3C9Y23tVUguia4FGJsBENUuWCY43kgFuIgMMe8E7l4R7IaVc7tdnE4v3gKOTDj
fkvYoVTTIVybl5PaPXy+iaS5IRaOvn/+QMFPRIZUGlSblSPuadC2b2PbodYfEF65sRyv7tPgV+V8
XxCZYgNisVn7GdHX8c0Vys0Kx3SPtEQqF4RVXX2tzGhi7pt5Edc58xYq4DhJps1/FOVqkW+zI4by
3Xrh67OX0VGN4GTqdwb1H28DyO3gprIQKJHzejbPnQH4YC5qYgKL7s6D4y6bhGx80GzaTihqPlnn
MtQsk7t+eb1HR9zStsNyRAcqp2wEUtCKcLeW1vowX7bAiRf8imc/2G30kfu52voTtBYeEruugsBu
cQHGos112xsro/za4YmrSgji3kwLv7KJF7M8Fjy5/CyXElzDsmuaAutTz29PjtnLyQubP5i/DPze
Lv8tz8tYOPgsEToDxe1YoCEzqJ9J277xJpH9VIe1VUuLJxEulEA+8G8nBjRvUSLqhUtgQ82+Qg9N
BcQqpkOmetb+m9T9s4IaxSTfWoFa85BAe/a35j0SWpdGE8VD5jEkxVZcKks1c9QUKj3S1jNrc1mL
3j9WGHop3792vQk40rEvm1zgA5lEk0mTj3GMyN6bkxDOENjiN4yBGoDcg4+Vo3c7yiu+0ZhGgn23
Hq3hozLkC4HzNhfniXTNKcfnYE6ewO/n8E2l/u1Gw2j0fHXOfvPBIuQf4JFvT7BHZtCQ68pMuWE2
R5y0e1ufzO5hs8M+s/ELGiA6unQR5TXayNqTqseEtQNofDrczjfXd1RO573PuhXXEnT2hv9YA1J9
TJBQRIz1fkt8KFj4BM8914kd1B0a9qmmPIvJa4GODusphrkEVjREjr/xSYoTVn6d5RNj3r59alex
Soa2mUcYn5qKIk3XZoq+80HJ2bIVLkLoijfq4ueoXZttRZEMkMti9tknK5yAR1L6sL9RQHFwjMjG
6sP9yaEWGAseMy09By265y85EmN6WtkOGXmREtvigmBAecUHrhxop3+Gy05Z07lkTtDPa9075cPk
EFzrRLWYsb3a7LxsuDxmTW3RKbAaLNEY4tTX0311ioTxu4EmPdh362jLeRQ1utjfEOPzHQOmXoiE
M/lds58nxbcnicLK2qqLKhHKgztqLGgcsBhlmFVQvSJM3F+MFZg693PjjHBKPrJNhUB1Zge0dZyh
O4KKTeVEju5sOCwElF1WwCGT5uZJXPpIDtSLfARxYxlu0Y2d5uP/2JXEHPNdfuCMID73Aqlnk5b4
ueQfvXI+6RIWm6iGXmHuiH7jF1C6L+eF9a7t0tkZZs24rsaskUaWcnR6CWUiRG4Wlz529s/gBvsY
aWUEpxVYwA32ebOafDT3fQPzOKwa+wi55zeHmE7VoWKscKwmKuf4SJOS9lJdRAWX8fofflpT8KK9
GOYW2xtPCthJOBbB0wX/w+XFP9qiM0hfcVYtFMQkRK5kpbo+TYjueWeVjpe65fa2l4mtD0m5trTA
0/8bkT5ay9y2MFDF8luWHMCqVdBzIyGacqMTsPThww/WZbJgbl26rj0MWw1Yl9dA6WZjqvfqLoFz
EeHFBr+lXSK+b5dbCd66qjP+5XyizSSyIj7krIXu4u2oNPwhY76uSvwrPmhjaNPrAcdMuUHVSJ43
Z0BoiYBnBM3mChhGsPR9DXcf17jT6M1Qz6tO3mkfYk+ddE9lymLgwU6/qcaSqWCWN9t0zc4ByhD7
gR0rOC+jR5oTx/RW2SPox7uF3TkFKQMIsha9lgRzQ6cnbmffepSmKookERATAYgKnI6SsAaUHDBW
ibdnaUOjm8nRUSd+KOhWCAr/eNI3+S9jzqhQkTYBi7PICfK0O1EJFrVWYWBcvLkX6zaGdvsPvXqW
AhpFQffqxatzPRm3XM4BYWAKUHkq/fzMw6SrvLZR990mjgNwDf7VYjjqyOwEmmMkVArVKXofPsWN
3MhVVDzzv0w7afq7Dr48Q+mtgZ4GITPBKPtU9klYqnxnUGpoK9DgJq3H9ug2SCxOXDiqTFu8I1RF
hmoPG+RLDtWOBebpr0TV9Rm+lv1hj927m+6f3wVyG4YREEllLcC0LtkhkENeLflxjh9l89WJnHCD
CSSQPhIuZjSc/pTTFjrLgknwRSIhOHzhn0YUiwwVBpWWMO6l7MrzIIXkiexsAMK0m2nvXmvCwjT2
5R6t3sJSOiNhFvMt7nI7I6hSm/Kji/Zk8OLYHztD62/3jtfqBSLAiq0FxsS1+mOfv1EvPJqAuupY
tSIyEyYn7S2U088+H85Z0jloMHD/2tDqcbWswQJtBfxJ3e8JZIfHS9GIt83zWmBHQd1p3u9npxGh
rHjeL9oqD+whvy90ax2I271s/4iOaGQtqcxILVCRRu7XSSOSwjlL+5DecuTcQ3+4nUr0+DK/NJf+
uf8ZNjt8Ckv04eGumdsCPHbNfOHOKuzNNAp5B9hOwNs/WPUB+H9S+wt5YNkbWuR2nUsCKqeq/nsU
1+B6YC0nGOwgVov6blIDGdq5H7wUrf8aeRT4pFdfR++D/z0yjacBm6+UCdo5snWXkhy6hrJhYYJB
odLWAbHEt6MBM3ehzVh01lI0Eintd7wMGRvDct+6rRkXDeDNUaqZrXPcRC3d7eHWfuR0CEgROpdt
52hoUM5OROwD0sirBKwvgewFK8HRIa7mweAgJhnp8guH9gxS+gCnG/SOxVLfFeO7Upj9VH78eNAk
DG9VU6Dg/PUNujViU9/+gqiew4deiXKI9jT3lO4th0m2tD3r1RB087Kl9jkQaKrw6yRRMl7fb9+F
S0iEAGEMF5r6bqWAGjXggdGIRhzCQm3HIvtotsB2vAAz+VPe727h+1MiMmnmxS9rfuQN867WAAnV
lCCi5SZD2iVvCFkLq9L6KiS1jfdWHX+IwGLXEcdLpvSLgfSYVwkljsoMtnIYvbl3edfxDBAXx/QQ
Bk0/Wq7Vm2e4AgT25TlRjW2ZPKwIV5Obdtso97VSg5x8j6ynb0AnUkvAdlPcipcIbHbWjNnQYG4M
iwfX/HSrDk9581zG+ipxeDe4zYYmFcA4t1a9H7wM2M62OTuYjE9dHxk7Fkr/oiWXLct8FnSYcow7
2mnHIBUKzi/gwWdAgSXFlZp3ENLhjeFGz4ucZc7p5ipXMCfpOxugDTidDx7eiJp2LxgzGBuDD/tm
KwbwaGa7M7q+m9qVtiN5RESy/JqUphSqxY9gQoGB8nbC5R22g1+8tWLUG9aGLPvDfrH5C8kea3WZ
eThY3VzVhDFyGPXU1E5CMIpYSNZ/W0v1YxFcFpmTs2W3CpuZisfJs9iMBTJ7rnOdkpaMqu2MsRdW
tr4BNVEpZaChP5VsyleulidS5GT1h+0MFcFGfTfMqspTPRM/CWpIzZGL1qxKMQVKMG96DRou6EtY
AeiJR0qmR7F6Dhjn36oaMbJ4tV6Q2DxA9L7sZr+ZQ4QJPd8KtOYI3NPedB+M/LGWeXF7C95aQXqu
UL+TpWBMP2UmXJ+b8eIkQ19IC4uYt7TC971JpZdbIoCAJkLYAXIZ4I2o+BEXgBcHqvA64/iO+Wr8
ZGtVjAV8ZDvVv8iw4166Rw2u0iQh4AwhK0kieJsc56uWc6hf4f4StI093FJXsH0qBcOieQXiYlrl
b4rCiU9UnTif0x4tP9SmEzhTD4NEvanRllNGW0yCI/hBMjMKZc0pfVqfW61asqSC4rY3jESfZURz
yjPy8d1pjHV2YeDUy3AE8Ei4jYMIRk43SEg6iZEcsnbB511dQ/z86t8F1SnmRapucmVZ4GA1+YEy
5m1YBwRu7fa5xI3Krdg2NKwq/nbgljXsgsj5bECNbsc6tGu6Je5+cuqf3TWoIpS+YFVSwgN4auIS
f9f5mVoslZT0LYC//YYNMezWOXOfgM2emScHCvYyxbWm5XCXVp7hh7RNovkfM3blEGUwsYkOgR8c
8IlnkzH50y589HZwhUs2AUaDFZQm2b98b0KnLzdl6XkgHW8/qPdA6+AMh0zfWGKBBLdo6YKdY70R
p66W71FuJ+n+tZm7IGKcQTgjN8gk3pNPY2AaT12R+CKo8+22arZcqqUc6WER01b0oIg30XoY/dUW
fwludu47m1Z9/4wHG1QecjlmcouhaA4XvR2/q4keuCERRJxFY5K6LdXmGyBKylcSN/0lr2FSv3DQ
B7I4x9IifD5vFitsKPGqwQyuHIltuSTqQQCZioaUecXcooPPtZtTGiBvNCcaLMa90DW/uOR3WzcA
pxmYVcRKBxevs+7+GhG5CD/ibdDE3Sh/OfsWi+y5FIA+ObfpicW0TuB7y0l2JaFPD+65joHp0bz5
iR5Yu5SY+z2ytLjyChRp3RKBUcHaD/iI7lYzfwcagWlejaOSQ4u1bsgWYUTlTZrrdiDglcLkihgT
XLwJMVbcAXv0QY0cxpTwa/ZV4bFQoRsi8JVSEcDlCqye52/PVhBBK0ZRPZnOLKNXzBrjQzS6bBNu
XOPVtlyDMqHP/QiSvv8jD5wtck0LQZY6eocDVRglZsyQjqRW/Pa0qHONUXm4judJsfB0B5a/Hm+d
DP+FtMI081C5go0BcorCLEnIHE9w/bKsTz09j4PQUjpmItduisYYhabB097UZ4WyRbc+90wchavw
eAj+inPcdXztcmefGzjskIZ8yWaiMgLORmpbIp/4PaMV2PA8bwBk44tqNXWO0khdFhjHCDG4EJ2m
R4Qzu7r/O7kHd2WVRokdCWlH7saKfahyaYSdHoHzshgIk5wA2T1zgXb4uuXSUeS3v2Z6v1/ZB5x4
3AZxs++p+lG37nwvvev3rBKr4se711HcAjmtVmtOH4n4nbIPt9mZEEUmMZ1Cl+6GMyR8T81VSPOq
WAkDH6IvfowjkYE4QX9NT5OkkTzQ8C1/WXMheBArp+Cyn1a3Oh+LxBz6xR9qE11LTafdj5242XRE
t/X4XeKEnmhQ3jTpx4Ebu8MOhODAqG/aYNHeKwh77Dt6Hc8iaJi2Su7PJKz3YbIh10xWTiAfG+89
33VCbLagsaB0ui14cNCZOHw3vFH0kKlnVp2aFTQV77sV5cmhJ9jZyKx0D5+b1IoTcEtHKcYm2WvB
rEpjHFSG9BlTUmSyCSY9KcjJ3ZkDlBR37mUAQxcBVGLAUEJEn3zy0DnJkbHqZlopJJRnVActZ7IE
hMj6pr+/JJrjUch4BnWotyS5m0LBjdJri1GS5W/IKUvlzMa2s85/Tsf9kCl3DNrmp7hVpYDCc9Nu
03FwfAwiAq3uVYNW/bvUkMZfk4IodYVPjzav2s6NXTPYq1M1aBdSNOCqo68A0qEGitVncmlUcJUx
tOOY/104wGCzodRotcfUxbrZnoKW42ejCJqI7gk47sNxsuY6ytAc1A7q0UxMG4uGWFXbra0FlhQ4
dLHfYRnlXo8lsf9l+Kk0VkC1qhLM4SIfJI7XX/BKtGepM6c/n8kTYqOOTeLx2x7M9BmpkaeTY5pd
cR7atd+f0T2uqUDTGW1/s9N4hxo0bO0FFfYnfK1u5q3iOXroIkljqBLvLaZiHOlJxukx0V+erpaB
f9fEwPBsqV3NCODbpo3Bgcm6TE0ZH6eNdJidTRTdtg3HLDdmmOV1pPa0RmAR3K2YruJiGktwZGlD
MjqI4UXKqDkZfXc5cqjkF7Kq57W/joVj2ZfM17gS+HVv/VeJlgj8u5k2P2B/tFQqVCL5pbqk1X2j
+ML34MDgO323rZLr9oXihSicoxQ8Is47mGjg3A5rp6kgE9IWl0Yq1Xlqp7YQNRfqH8CGrsBEtB8f
f81874jLyILAuFG8U+ZcIStieyVOKr/BdJ69PKVGcT1J9zEnO3AVn8z5RwxMe3seeqMABiHHiTSz
f8qmKzrloeuVsYoQEgofd2sytfwUJCIdSR0bhijY8kKAPj6BIjZyaKQOS7Puta62lOeH9fPi13LE
23ufifbcuSB6nMFeFrlAgtos+CVAAKPjzV021570zi3AuMJp33YGK9U9m0YnqW+QqJAMO6+mTK3C
ln0LSea3j2+bf6j9A7AokrPnNCxO6QWylCVLPwwomZD81jAmT+MGpG18kZno+Zbcw9CUFQkw3/OW
C/TYTSpMhD4yiS6y2sjb695XRnD30IoyWkhur6R0aPtaSuBAPsLk8B4eSG8u3jxRvoZfODqPVXeZ
JeGugVYG7/IVT3oXBff7dnbIMXOgQabYFry+21SDgWOzqlOjgwP/emLZcT8OAJKIH5110+/0mGUh
N1ubKjW/Z+NQvtiLnXznoPnxqyUAwll2bAhbBlq72Opu7/W/xUAduJt/hyHEwXbio0optNXMp07u
lRwnP2mj1E3PB747JPsZZhQO1o3q4UYX43DRgISDz4Mfi9sGNDUvct7mMPEB4hyJl2+lyaurFLL1
H4PYNzC4QpAMzCNUejqi2Kc3s86RLPwWaUcwECBQ6EnMleKMc1NBMySRps784phdhEUUho5cUF/E
JNcpw7cvtWq+O0IOFPLXiXt5QM5asGcdhsPF2oo9hYAIzA2UnZSXBo8qzSzYuqnF6x8bZToauFll
xOWhXiXtNTrRK7q3kYff48gBZY921TMYSVGmVPIcw25fDmbi+eVwF1qeKhWN0wey5QkzxkkcsxY9
eeVRpKj/EKCENW/F0Rc5+zDvWK1DR51QpsM+vd1cFSLf6UsV1QMYI5b2UnLpD+iDko303MuM1k/N
jz6irnhpYkKvjM8h89plNhkvmA+7snme74z7g33LZhpaRKSqFVQKwtbN4iiOlDUmmwaQI0n3TQh4
8Hp36Y8Up/sSHbQZO50DouEVmnmFPB5+KA4acFmaC09oeot30XgpE6W47N1k3+sVwNP8zFG1DoU8
6FU4FZYjsVfU9vSn2i4wpBhFrSMp1pPwO69eqQZvWN3CAp1k4wsL8gt30HSXvkFaNjTfWYwWd9ae
9muZbxQ+aDyAB/iTmHRI67DVBiGbJI+fwHV+LDyi+VBzD6g4SxW+KdI4O0r3aLYQGuR+LnnT4BFs
GhpOiCd3epiWhEBh4cUhzFlaOWdeR0lMcPSHoWXFktUr0oqszcS1T3yIUNrObgFRweJ4QmUvMO+6
1J+mz6wZPYtkucf0BgsH/56l13DMTa4+b6J1RNJaahVzX8tEDYzean0d7US/Aig03U8r9/8dmUGx
oK7XXVq2bIq0QC7nF+7O5oRHokj4M9Nu/sQWCKOnZ74HhcEkHXQw8AC5q/xEtBFup0qpeMeDiRDa
mmW6lIygECT8gcSAJmd1N1mQRBztEjlF4LljyPq2qyoBN5spZQhaH53e/E0MW2T5p0/tvLlaw0Fy
cRBlQxRrVq5asaTruExI04/ZDMrCs2s8lLErn1gXuRf6V96ydTU/106afbzQt/HPtd7Pu7TmxE3b
co5E4OGGMidB9gDM21AE9NgPJ4qdgj8vcJEeEGdGh8h+fO3NShdnojuo5BdaBk++ufQ91lZZsypy
GbZJ/ZnMeEze8waM6bDkCq9RD40xKsD53YmkGA/9b5BZZvCniw26ShOhOrmfGJP4nRMeKDR0y5Jm
9q6mtvsYFj94laLhfEvwD/dOUkEo2ENyQkQWNDyzwnfQB176hc4THeEwnZr+jnu8bB6dXu5gn3Wl
joqbfJBqIVhlRbjxws1dSi5xluPI+TDTYHxzBA374tn2eZHy+a/zoybjZSQFF42kBEuuKDtxeugP
tw+lMQDKPLMLSfLFMt+R9jnu4mSo13a7kq+pPARyO+H08+oN9d90ce36iC6tFsfRrziw3QS7hEcq
l6I5pg3cwWBHwxMcq1IUd6Udj5xxyOWnBLFxeLu/0mWUNu6Ev5lc3ZCA2ULWTGad6C28pcm7kDkZ
6TXCoz27uoy/VgxuKTYbePGwkvPbA6q1NeJ8qzOnqs+lxCZQjOTjcL54wM2+ITXSs7AFxVeLvzsv
mdTvMTOFBetyUgOydhE+6O+LlbOuvLJwaHHoESu+xCkwhUYAAdPKLxhBSi3cmf3HJa9w50jBS4yn
hX26jq6roWGXvttHQDYWyZxV+i/93/PMXAKWJcmrxmsT5LIB+ZuPmVyQ5rjF/vqJXQTqGrvuM07h
HpH5B4AZ+O0IkkAXY88X580IDneLy8msjnEn/4s/lAokUhTCPE5kNGaFpLyy3w8Hn055DKbr2nTc
TWFaCQ8sHwkoSlMJE5HjdUuL70edVl04AG09LjFRQpzSgNj1udSLtRBuzDFKMiRmN52IV0tBpyQ5
84J9PTD7bVaEu5D+Z+/k0WeBgY9S9NT+iSEs7i9IhF9HYdAPqmKjVWGXOgsd+tjlU5o9lPgXaNfy
IHrrbuxcjY0hmh7n3cp/dOh+3tiD3S7Z03AqMbc3DB5xaRXL/1m3OloKOMKae62cSnl02tX+bM4D
YCJTQX06+zwIva/pQZsXHlfMl/3XE/K6aGDzkiT9DgTm9kMsoY2SzwtfT2BRCGqEilwWBGFbAAUl
7edrSTnYTIk9DcVrgn33bmkRumblxqAMtkgJzQTE+3rxs1sDX3yLYuw0PxeCeSJV3g0RL5YK7knS
ZA0Lx1cpaQfeiC1JfePmGMrugi1NEgqhUtJU8KXSG7c0Cs5bRZ+q0mslNNqycExGYG4SbsU+GjO5
skktInYDNBlAt53GwkfSS7F10stpxgGmETojxYS4LkUk+xdNln6r4wypZDB29ZbpDXxoBN+NOaqJ
0JebGd0y8ZXa45TZaFmXQQ9cVjvhuBpTLDJ0mWAzTEY9XJ9HjfOq3J1RfLBgztlBF6zNW/Kffn6T
Psm8QrB1BxVp7yOUCOaDKyBbZN5G6Kgqe+GJdCgsuFqqKK7aciANWIoLM3swDyjq1VHKxGJ7NI+O
eZu1XYssOYhnSfX1QzsxLlIp0ti8We2Eri+g6MRlJ49fpkKuixFucQE/yaAaqul163zrFnIq1Amy
KmGtM/DqxbsIQlGZyQmes0fNO45wDJmDW5NViYt6EPxsU9smleNrLCYz+hG86Z8XHOrdFH8fr/hb
F609K0/t6BLtTAhS1w+wPIWWoiUuj/GCGN5dLd5QJPatNs1jnB6ieZs3CZV4v8cS6K78ra1CzhMx
cy6rQh+qqxIYxrs/VX76yIlbuWlgBX/Z8Ph7Q/WqADzy8wlIjBSnp+8HhI6LvVCrglZyYE56ksVd
nnMRm4HZq7VvqYvyztYGr9ZI1V72emX2mW3mvdgCjjwVVL7GlG7VjV0jkNj9YUSb+zctuQo65A5y
TkoT/9eoGBssPSSv8i0KOFb10YR/Xce/Nl5maErY3G0cQMhgjmh29KqahBz49qJWc/M/sWuO+mUO
7H4KhQgsFkQNaCX13P1HKfp/m2Dp+E67nQijgM7OXTrO3wcX9jnULezsxJnL3S2s3RLvqGQKxade
0SFJO7LjQXPNuVSTnsavWkcysG1uueiwo3cvd6NjSlqIsP4eLINVsnfivwcZk8gytOlmCu6dqleX
T6/V8XzNYHMur5HJpi79+8EyNToMTOo7upjADtN9i2VvL8qGqRzKIQtJSTEVEuT9lxz8f20zb6eQ
hAoeyeCwF1gdvfoWVqj2Bq8o19ZqbI2V1KPppIXtnZJuQSDOAC9vYY5i/SSymu4ZyR09EIWLJvwv
QjH8LX+O+TVzkTBmdCeDK4CBDcDA1Ug6enFY6iKp4hwS1PczvoXKAf3IRXBBYNgt1I+O8HF4l+3d
OmFY2jR/2VjpiJlCMosYGlqw1E2rQgEsfsnJtG1I7IqN4RGxIja3zmUzU8zAS3ab9WNWnbm9eLxK
gll+tI28PzKsxyFxa0yCkfshUll2lEfQrRElToVvOZcbH13bcM0W3fyNmdio4tTm171sXmkHVRmS
VUs8DCU0Wcq4z30h4IWr5dQTYjw/d7SYdV6M1hBBpWCDVwI5R7BJUpVZbSNDUQkNvBlEO9r/VP/l
3tx1yNox1CHRyySTt9su7Z7imEhSKdUuQbYnDHbjjpYXPoELaJJxewVR1WZPfluIdVWjHi0XhrWS
ZhqLOLUTEU7ehmR7LLZkLv5hmRWt0A6nAUwC+wphEw6n8y5gnl7hsa06h5UoPQ3L8P2VO8CI1jUQ
TsZ2w6N3SrGnn/u7rOrIwIAEXULCBsQYKYEaBrTuOqGOhEmSCDjEk7RG0B/UlaRopiB54mAAMkl9
S8drshjREytDTiB5w3SREJMUXuKefY1h2bGHTp2t6aypUQzQQjSKatJb7u3vkSndzU/MSN2ouvls
5JQC76nQsmTaAkWmnG/H3UyRwAvFjlQi6H9s50THmPYsRY6QuPorEeptsmVdiqMyzD8lCTDcad9h
oyqNbTMuItME25J6EveJlqwnXxj9Yryb3fLJOSX4I9V9Be7bVquz2FxQB4qwN6sINdxkaZNHTYw3
TNCglBZqVQ3FLh782PJC7kOcVZugYNWbtd2UjybpcOE3y0lzOM5+RrVYKhOVkCXo0YqNYNmdKrGE
3vI704fsVJDKyJYu6HExy354XEjm9HNmuGhR7hvUhHlvDZGDso8nUju7IFIovcpIHpMe6568Fp4F
JW5zw3DmYwrIbbuysXURmzoktcLz2CugNKR40u+pFq8KlVPiPDpUMkSwc3ayPWA3e6rwk6DkGU/F
ZnDxgb6Vu8LgSlStX02iKMA3YnaY1Oogk3KVd2McDTgiuPCyELzY0f6gokjNrWWakAq549CJmCj1
93fFicS9BioI4MRMAFJ4Zpd9XCt0VF36uVKHgchESb8qO91PLW68JevRdYS/87Rq3FGE5pUrV5me
b3nEwFVl0LnNz2a1w8cLN9fuwSJZjIPfdPGHYawXlIwRUhPUvqRMjRi9hMsCb+bE80Vl4c05pj+U
58ICKrM9+1e+WGqNfnPHmFMfIuUIRB9O+PftUqsmgTNlOl35f2zhnlPqjqkpxh4R0+gO19Rl060V
qpE8tAngAI0LPN+JMqqFbbXM/IXYFtm9U7VG/gN7NlRGzDVfQB0vYheY4lWVv/FGSvxUGn7z3Jel
SXo51IBmNVMnUo742O2ILJicRGBp7BQwmHZDqANV4fxMSNU+ji289WRpwxbfqnNivcDWc3klgulB
ht1XqhASGFkVOzEIDMqU1FABg+svwgyokD/dCona3UAx8Ma66bA0rDHOWxXbvaFeiGpN22pHRCYh
/fqr8+73dIXHdsC7rLpiTtEXh9iRodmPsrWUqxLvzvi3BTe1W9xnKgFjeWcfJAluFozPRqQ6SITL
EpYYrTu4CdGdLO82yqpjctNcb7flY5hYmF0udtWtE9LXyXEvXjk0F5GwHde8TR16OvxADPqgkK+F
83xtnkW04MLzLbhf+fvlKgv/ch9tqkcnD3bFSf/t8U4X0Lw3b1Dv/rT1OclNWuOECLctacpAlg6a
pIaPmxCcVYWqt4Ceg9JFTMIl0KoSBhmzGDUSjEdeAVOLYM4eVcSKtTfJYb4G6/PySjmSvrLzafxJ
hJxorIJ+yTDT5mT4LDJYcP/hMc+gcmukDBmeKi5p8Egm8kZbsUprFvHvF/q4G4i18sWbQVz8GgFq
GmV+ex/vv5thKJCW8bsJI62kZ2pNMEYvIdjQuaJZpDK5TfihtrQegQdTvWotkgT/+wVCQU5QKsah
xEOL4n5ngNMfQl/l7Ivkyk+dnskAVhzob1+FR4BX1NEooKEp2mYuM8xuE26x9F6m8ADRNsUYRW8A
SNkbSIW9ulkWBOK1eTkD7v5mqESS+uw5zPbdyPZc7mjOMmZE+ZNRo6GooscyM1KOvu3QZxTSIGCZ
MlyAmlNR0Snewv/XZQAmKqeyPVtZFkRPzrLzg18yJ8jVa/ET9A2YNC4j0R9VBM584m6iEYhd/RCM
/QleRwheXrjPIWd+NLSJXOZ+T2G+B83BqwCpCVNfhEl+wXtZI6lfsbql3OKnS/RrNQQ0xsQexJSR
k3eLEBEJ80Aeagc4bKdlahaX//97APFrd2r+Aam74lQX3igpuB0fO3GiIKugcversdkOXdVaGIQy
b3bNcDSQKU9QgQtyBq+rcpnHJ3kztksuG5/F3PGdCSB1vHX56FNF1EYtNK/jKLDNn2e9FmQWnKKU
djdYoaFSqP+iXdvv73SXcXjhBVR3D/2vbR6M3Ys0+DeLW5HbWcJoRK/bolbQTXdVUkxaUOF2anFg
qfzUwu1WdDYRNzAZWRlCwHNET24Ia/+8e8+0QmYI/hwordrEzgStG1IyRuBvVebL4GKeUQ7NfNu1
7h4363ubJGEs+jDNMofl5e+PV1HYV7bj53KKNKnAcnS45sIXRdeiOXHnr7mz4k5ZT0GgcxaFcDHK
gT4o2+w8SZ8dY4kUPMJGGDSJwic8x7DrFbBptIDLGIbJxu74tIIliQqJ47Nzfo4ql7WAron2CKbX
MhE1GZ0hdW0tmOuBbOlC0/TM3tXfz1xRNuC4I2wsOgja7kmlX54+PoguU3o6IKuuNW7VFxcq3DCU
Mx7drRRE+Gmj1G9KmQXqsZyS6DsONTZeE+fYNzr+QS/LdE/YrJdLAiQsRD4BxvzmSX4kiiOg6pjF
OvxnVDB1n0nGcz2Ut12BND9t4DUIpHWxQeqZ6lWves6taOraMM5u/g+qoEncHID8nlny7bvyvWsU
dQCztkeOrweyWrwQBUXI5gV9bVQH3Q3vTxeUn5PsuNGnrmiXjsL/KbVpMmo5fucya79y8V0Tzxqd
sm0R2kC6ZDaVRjcMNyQv6H4xRaOnYJyt3O2x7GGlzJLM+3XMa9V1VWTDHg0o9IT56lMeJ0UMBRVu
ayvl4nx9Hlbe48/kOrlg2o2oleYYB1KzhiZYrr98tTgJLDMCDoPTaA4GYaL3RpLNNLyWF1KccMnq
HopI4vmMYRmemD2LKkbwn7p3SWKp3KgIwnPfajRTpy7OD/7RbKFIrUA3TjyhtYI+yDIflKpxfXPM
/Dns8Du/0+s4zr7Jo74FOy55tWFkWTelZVhTjcp3ZU/m5rU7gk1FZNg5DUgxl+QKvC942MbTkuwS
EAUm1UohocPm8vkD8ta3A7drwYJCaQ3G1k0EjfcXtj8UlBTP+X61XtiX4GkREhVKqNE/MjBWlSQ/
/RI7O2XXNoGUAkgk70HZ3SkMKrGIHKjbY1ViHrN2yy5l+SyQwfywTzaIsECUH2lpVNo3xdjzaG8a
aMLbmuf2w+o5RsPLIP0YaolUy+Xtos3mb9qUaoedIuTCyvbCu8fhw+rK/ML9iCpt2a8Pc0+Fv4Ff
MvsS+XWcNDQe/4M8Vvue/bZACp1zFl73e/nwQI+pFjAC6Hok3GRHb7L/NMd5Egabfmu+7Oa4L4X8
DIOraXhZr6eLHVLFdi2V6NFPTM8ciuKRzIVA8K64sm+omboGSpPPLVlcns6v3b4Il3QK03JKMTDe
WbOqrURMGSXPJda+vTiL3cLNgNuaDCmvPeOYggp75Fhk/5zE/nW0tidNTuZBBZ/gYpCaRL+Yl0QU
UCL40h1Ap/bARFeKTRQmd2y7V2QWKx3+w8beM6g1Py6nqU1FbCPWEtyf6fAQHvAsU01cvrIMR0y3
nFLQqSo+8AxcS+6LFu/vSuP2V8OwgCo1FWH5uSRVYlr1bWVYbk1ou098pziaC2b/wl5oHU72jB47
LSk+jGeE11ldln0ve3kw0uRJ8MBJAgajnt8mFh4+s7qV5vSKioB5/CV8ZLfH4eTnSZcsmnhjcawM
4p30+bXes8PNFanJXAVnOtkQmdSbETT5H8AYVmzdSLf/CkHzJkBuxntRtDtPOoxLQ42QsFzPCxl/
AzazXshgAfoP5amRPkvXNNqNVM3llz2OJm2OD9zpWCEeqdM+siJ12JRi522DaQY46gEg1k42B9+1
igcccBz7+kTqh7t0plsonwSLpfdn/KD/hVCOVssgTfoFMkAOBMoStoKVocdUHsti1XMpL8xHYaT9
HIzqNRzrP0awZ3Ct6p027ui1c3bx3Fi0SXXSJ/r9k2uszphrv5PATq1G0HSDgjPZRC54OV0bpQiY
uBIKvzu8kZHMNV8riz6E9uh+uvSSTzgvxnl2e2x1s1a0mPZZdA7yTffBU0HHjjNav9njjU5FlYq6
Tj2TuPUesmLiElULfbSCBiO7iPqgCDTk1zfO6/5yRZRPp5CoYHdsE8w2uUhqDu30SdFg7z694cO5
QuFoW6KFKdQo2a+pfMpenNdQcyz6g97LAoNbkymvilql9u4RDBUYPvkQ2ThQFYwMB1pOb/DsiLsk
EBY+ZR4ZDh2/XO1ZLc83kPabFf9eIUU+CgmP3BYP4Myr9u6ElEk1VMSzFbjHR7T4+0Q1ycyfcHAa
RoNeIwiq+9vmTzYaNAkv+CIku5cREiMYL92hy78j5dj3F75flfC12cMtUNGX1H6ALzKn2X4sbMbR
9npFdj3ScZVOA9nz28fpmJU3ouAwTybcLyDYxStl4VwiJxikW0fE+1eGtpdBJrApooCVpWI2ffIR
j5x/sFgbUnmk21YJJtCBnhl1RFDYTmlQc2hqJ7HNMKBJ/5axWUMAp8APVxXxfDdLx0IMksXYZPo5
bfQA9R46KPgrw9bVeQE9gSmuXh8WkusQw8YkBZMA87hphC3HAQN6erSRWeenBhsG3468qpqGL4gT
Oenem8W1DW/tRTa0M3KCo1ssWtqQhfqCQL4Y4lxM7Tl37PLtuIquXr0SOOv0vENh60ONrRY9c+tC
uxAOmQ7YxoSRsR2nT1BY2pOjDi2RyURBIz2AYDaBiHJtFa3oa8C+OavrKy02LvLIpNX5waQue0Fw
lis6kcf2HStz/El5QpgxtslGp6mF9g6LB57yybo/uo5sm7RbR2glkKYZgJ9684JjKNTOlAfnuDzF
MrJmJnMqHGE8EeaH3/L38Bjn3XlOnEIy+in46uYgVPq0jSXpDY94KNMsWIcn5pGwlm7Z/PuM5WkO
OnXetRvCD5Z1Gwuj+0+xqCS8Upucoh5OgullgSGLSBbKCRP89EHv6IjeHw68ImG9EOBInFpDHnD4
YM2HMGjujwVboZg/w4exYvzFqmDWafOHCbqMZjlY6nASiqsPvhTJrTNZyANCu5b8BY+BbfzHi+Qw
m5Jp/Jf0cF4UpdoO2OTuNm2px4CB6Fhiqiia7kO+LnAoya5mmITTinrz9sAj9Q18+A7lwRmAhUDx
4fBCJVu+ZYrYi+2QURrjOnXzzYNpCvGp5AEwhnNnyBjOz540Spg8LO6zrW3tvCIevq9KFAPZcCfW
1mFCCz9HxNFEijTq8DydAkiRhiNsZ/TeTFMMSus/I3hUmCtbOfK8173F8vQPFwStNQN/Czo+KHzO
XVhuBwL6KR9oPUcoJSlcHVTA/4B7XrLU5VQFEqDUBouKC8Pxpg8iOuR+V843Wtejy5QJpEB5xCWY
cwrGQHBrA0m9DlkCqMPck+zyQ9L8JgEeECZlRrGxrYdmRqYYYm6S11wwfLEWomYr9AQudrgzhM9f
cYgPF+77A0PUyctP8pDQIampYeqDnwSInWOVq4GKzWKciPPbX3a4q/x9BSBafFstwPni7atH0aBx
GNgRvYCiIK98GFstIRqvuPZ07h23xca73uG6JkzenSDoAfxzB9VGAbhygNYlNkOCZ7srVCS1DsEK
A1mao6pz2srmBWSoW2UtYIQUs0g2DKxlaWrWSktMryID46+W4YXwMokPHv4eX8Pw1uMuXDwZJbvp
s+6N9MFccLqGKx0uuN/9HhfE9pr44fswxcMvijOPtMxd4lVBJjQ0WT2KsCmoKYUTuyhIK4gXjBM9
NMWBPRfa16krWxtRHRWR/8vHgXNvd1QyRD7CAra31D7xyKFvqnrsLgZHruQ6kLIBnp+Ii6PZb4en
3NgXftGb55LWfDNJMZkOpw/lhaVAxiy4i1rW1QCH3K6YCLaGlJeZ+qZ8eOI3M6fSZINtwF9bB7G/
kRKWCYkl8sit8Wod8mSjrk6W+ZauqPuXandhi+yIq5KsP8Ig/SKfIrshzaX0GQw0J8GxumUWH9me
PylB1Av4kWekXJe39N2osO2R2sAiOsalsHa86VXp7nN1Uc/i/wSax2WQ2m5nVPDjjmt5OmUzsO2s
j7mV5iV+i5B8dXtN2e0FJoAtUUao4j+NVDL7ncsNcrm+e7G35zS2T/TNW4AY16GnK78rYcXbJb1Y
pESGI0UalTjJCBQanCKmDSsoD02hJhPsxVFwqzvUL8rkNxeCxTjKxOmhpAHZEsniH9A0HVl22aU4
1oW7vrxV321+qrvkGcy7hDpQmBzwn0PwLjs+Zt7UT5tAgOx7sFM+aIzuAtRnEqqhux8PcQK6FYD3
YJV41/E5kt3qxd+4uVS7h1DrlVbGxwYCsHqN0SCBtG+Yn1V6gfhAxkmtvNLSj+JIIxawzb8Se8mX
4zShbRUJrAjvr//HKdSpjwE7xr4e7DfSIwao8h4ytZb/tM/YyzxXnT4+PH68r9RX1QZ9derffp3v
h66ZAzRf0IMo2JeBZe2pEXfgpL+VXVde4voXXXWeOVl2mJ0RI29yWnobSAyjk5MPgwx40RxECBSX
1W1dl41EWjLSwfl0TxL03wWqm6v5JBQZq0Og+c6esD3YT9VCpoSSTlMHDkxhSJgTsGx8aDx5d/U6
95jC9NW+R2ERtx4Z9E+23eSAYqnt/DkHdxidp0b0nTnO8cy7RGPfE4SZZ9BphxK1aIzED9XsP1U/
asbSCVF2ChAotmzVcwCSCoVOqnE340JTU43CW/IZMuxcANoqqC+cboxqlPG7IdNkiFWNEqioEvZc
GcauDNyUXj0BPln67YAeSqOFSzWKfFU36H0WZMCMzeRkspVMR2XaoAzMJHC/svX+Rk2sNO+f+2e+
KaBqitAyCU5O8ZE2Uxioe6WE9B2bEz3FiyPeoW1pCv4CIgpZaeX0WNC7bCv9dmPORzNt0R6ZXVkH
cogn1YDkCOMD5n+gs9uCBiFyvCwCvuiLMXx6wP/mcxVKErE5qjSooUH+vk6VB21UKCNToINDncdF
0r4kg5sJBrPuUy2e82uoQ6Y3T5yVQtzDozXPPAvokmqbPtGQa52MuQJPI3TyYXCMitWqiD2JM5Sv
+zfZL4DxgMricSIBFomhl8cnRRrzRpclz+BaG+PK4mg11+FO9QKgpUMQeQcRlj8vxPiUgqUyIvim
CWHUACziQlVM8NL3J1iQWUFr0Z4A2S4dxBGbY7y05uSRfBUHOiLKyZst1PD0qUfDZieVrHDQR2kE
1LDKgqNasvoj1smb8qOzqsWNM+6uinp9srVe3jp7gdl1uoV8l362rTrcOoYe63q4D/zwa8ZFla9d
czSM8tgiAga6paqcDpgps4B9ZPL8Qeu8EE1gIPykpKHecL/MAc2SiYRMt0rb+fnJ29mnAF9H9tzU
c3UG9y44TCWajvQZBpZbjtJNCU02Udx/IkX7z32AZ+TPX7KtfizMyO8TEub/a34SGxxR0ZFFEVyV
giw1/hclAEknllUjsQHZeRIHZuacuf5Jog+d19MZA+z7qcC/I3OgQV5IlKoQyeS0tpLpsyHRToCe
rzFjZn9+kqLygSY4TxAawZScSc8J7Ynbn6DP6qyuZ7hEhOxBMj/qrKpkeeXbth9W8HXw/BhzMO0e
itGl3XsZvOk6p/HfcrexgGwNcFyuZOfZN41KNkHzvi2GTeBIzH3Sz0U7MrWh2IdoODQ1MPNNAH+k
VlxJ1MGHvvwd1cEcI4y4hE361n++qP4x4O5t81VIB6cQy0/JFQrNSnoMNzeWbOIZt96RNVABUGzn
jZLXC/PlFmhaSXJbNOzKmKyN8YbflaTSb7/sS6GwL4S8Yg8RZwD9o1yBJQMHb3cC2vaBnEFCrAxh
FceqbGPXO17ELHuOlJ8fHac4muFLOv4b8WvG07dBsCu5TyvUK0oomDECroiOsn56ijkE+s205lJx
IDzJZP17cKQNEDip35/f7ga85CXoxRskSRaCXMFOzegmbxSKCb+ozn4D6HJdq+Z1C4zj10z12mmn
anbEKaWM2j0WNemAnHiyQbIWLKMuRoBDwCk6SP+8T4yuL9K8ZephjWFoMN/oGuA1IkeW6pFxnEq5
HnTOhhC7p3KAgpUcIMi8UFOq59ZlV89JeBPY/eTmsWqS7NxN2owtTVxoA+COuRRaI/lD1Svf+plP
gycc7CuSR1ixqHG+WmbsrMA207J5ILVI8LvLDRLYA5PvXCjjFpYwQp3rd3D/Gt9tJj1gy9o8Hwub
CFmJIhe+XwFEB23sYIysny8h5lvtou194LOutAd82k30xYCtf+Ahdc8twEpo5SGofxXp/mYJIlrN
fpf7TZ2C5+d5fBTXUWc9WtLTH3n9rNvyRL92kMQt/E4uJGsgkETj5rfiUU73QyYqMSJBR/ASBlcm
Ik1JtqLkTV8jFxJFxfZp/aI7AzPKWxAwAZpqRsEKa7hmfnPrAGjIj9wzdDKlizLgyBVr+nQj/CY8
2PUsDjexpFv9nqB4+z9FTN31P2S5FQiXhQZ9hzoNq6pw2tGlRm8jsTDExdFZ6jNI85JvAkPzRtH3
tzSWpApXaPz6vTGDCDhv5Eib02QBKGoGoa+y0AXVD47xJlI9PgJuJF44IllY+1VQn5zx5JE/4iE8
k2qq1oIlvqjpe4zyGn/oMhT8H+5EnNafbU3X3lznZNvd15nRmIBSpTMfFccKf454KeDxvlhV6hEE
zikljnTWRw0evpmd3ZLUFgzPQR15G/D9EoZnEhrhohrNT+/gAPNjx6XBmau7gNt7Ky7EoFiIXCLQ
gom1nTkOcCb5jtARHhqMlWbjBa+ToFJMmrAljcMikshdWc8xqzQ+uDY75NTnbU3nVeibxRpePYnl
jquWCsl6qG0+41uYSADgw/4jUWrnvIO992yo3wZWLBThdL+7FWcwhoDgHnWrhIv2EaBVzw1d67g2
dnuFfNvOsvoy/3idruIiqZiO7SqTKXi4ghxBcrEDotwzhLGJScJe5JOIUzooPjgx8kiul0/rWzC2
Hrt4JzlU9lVi267kPADXpqd77nVWECXxkh11QF/TH9Re5USoMf7jveUrVqGp7Fvg+VJ5oHJOl4D+
hHRwi+7gEeYBcHE5iE2gbUBqS68kDefcPb1kgpF87zlZ1kNifilaa76soQRngIa/hx0uUMB+l/3j
auAh46RktT4tIjPsb/eAkt9ptXvdDDk0G2vU4yEQXdwnXdzAO1PzXJMLqCbakzb1qyce5XDBBfgx
b4q2w5yxnCmXu4nHuMqHk3b0p4GJaA7ld7/WoCeQJJ+rGdPOUYbWb73UO3dyhvxGkIAjMv9znHjU
VAIZ1oB85vZ2U0aHMxnCfb/X+axDkP1vLAIHcUziIZQIGITN7goOifAGyWJa8VnzQQWRmed1RWG4
nwhSDFaB4OEqVGUSH2FtBl35uozntJSi6nKAsZxD4FeiVQc+HLsAdqYehfNtWz2Sfw9gBfsPCzHr
aP1sPWOgyAejhSUWFU0GSrQMQrCOFvIO2VZpsF4uZhLBGVvwO6xzcAmRjhnE7I4/5dKsasD1aDkM
/c+cb1mQKhau7jlcSI0kV8BflOcWepMJ+c3Vv9KfhmshMUrUK3gw3ANJCvZbOcPm/E0EZ9wHyCuj
6cgZp+cDs9o42taKDtFDzPTOfwyci12p8gNsKWwjMWP5IOph5wR5rj17CHNd2j1LK2XARTmk9o7d
asK+tfkN/CjU/d1iusx2hPzsSEdVcV8GHbQ1XqGEUk2BpeCaW39ZCQuLCACEbBghUX5De50iuC0H
iOa/OR3/5A85tErF8oI5iCVSQ8Lgrk+6AFKJdw/ZgHlVMThIcrIPlIhzCh/pGFaSzrriSHbiESvq
/4GCp3x7sowKOc/NUgrjWrsaFNrL7IrmgWYkwr/trirDXOhzDsp0ihgxojuhWtaFRVmPGDJ3q1sh
LnbFD3Z2he/DWH7WEh6zsDS6xKLWHqIk1bg+q0DkS9ALK3BGael9MMaLQbjt0/NVUFsxRQ3GaFxd
NeNvVmg1N0h1VJCi0mm6d+khOZWQhO55RD+vW1xngCGyJLKiAUNOiAz/0lJNG294phgr2L6HhzH/
VKWs5eF/LwOiOKmA1i2Wttyz3/aiRNRczQqwF8m6i+9Mus4C3UzLSqaAxQceVkOI/BtJmvwsab3P
YWs77pzr8P5/7GErIqWWJ0Qrxpz+AuXrWoJmJzWgTd4CgaZreQQco6xMTVs/+tsfuMwZQZZx3E79
PgnzWCObjm36Uoq+iKRyx0Oi6gJ2ma5Ho/X1br/ELg3kM8Gzl1v9OOj2SmgzNcJZrXkDb3sIweAX
cvDHb5GKVKqEI6hxU/mi+1LvOGipxUFyzhZsCubSUzcG+XkGIrddL8CBaeGgiSPW1XbldZvyYM46
Ph40WOOYul18hMsweV8ulg6+5cn4SLsvIpSRhSAMM0SSWrHSGBGHqUiS1gUSKSbGSbR5unkzH8jJ
WwRVfb2lYroI2IwCR8txQjjNgbwDhIH5nB4KwdePGjhzgMkcHbCBPof9FaBrhOk83TsUhiSd13OF
/TkjpMfjj1oFGWB2N/MCCwogj38X34KZ1dD4z3LjUFllNNj86e8g2nBTbRYzRkmgtSWvebvtvp8D
OOwFav7sZH0HO1mvxr4Ojum7aadLM7PXy5eNYmVwnStZzLoah2wml8rex/+zc6cXb+pVAPKGW58z
dCi9/amQ9AkIXD/WRi5rvxOer6crM1Qd2v+4msgxrNs74PQBv5EaKNmXcMpo4pOEXoMwFewjgHhd
E5mcotVwwk6aq2HClRFcAio3eQNwmwavcxTJn7m2sOPXnKj37n1vidNEYtDr8pZG05bT8f/xUmjh
c/n0brdtgwSchpVImU254EQGtRYJtyyOGssXeTkA4tu/tulCIM8UTeAi+rztjEmzAtOh25MIoh7q
CncRE7evSxPjC6C2OHC27/rHiRtgaC25eDZpvtphyZbVMsOoFG3OoYE+mJBswYuPADpdM4CC8fDQ
Q2s/5FD5BTUcp7FvaVT7DUM2thVf0bGroKlY/qOknZcSftkdMVFsFupxZK3MJqQyN2gLJZorqtNn
Z1qhqwd4/1jKDttlcwKG56ABfh7BOTcvPYgxsrh6yOVjkzFX0SSqX7wVpB+E7ZXkEXylFhm3F+7l
/3io5KKDoMXgvC6q9OGjXvxoXHJqrpbOwcvFLF/4HQIt7wRlKHvB+TJUi654S07XHxVIjEn+HvTF
KiZnCKQGJt8PimqK1nCbfXLBdaxJuVwtYLPdpeOUy+XI0N1MOGjB7L8KY/NbMFmT4rql1Ybob1DB
NWyd/OjbKqJ5q5x1jz0oOjb349KJz489vC16u32XITTqU8AP3Us5xvQEwThgvls9UZiqZNx0K5CI
ehrX8P3XSorJW1ZGhD72ieWqTwAmLpUiPCktPVVlxrVianW6deNyK47X8QCzGdEUVOS168EVm3Ta
oMacl+BmLPEGbxEn3b8Y+MFJqFZsGjDf9UtWKf7n3aeyRXO5C6jqgKy1qUDCuEtugurA+sYi7IdO
yuJglD6RezJjOnwXLlz5mENfR7wbQyQgnTOMgtx1Li8aLPzLOGsPq35U8QMB7r7HR57zCXqe/PdF
e4oOMAKy+edh+lQyjP55Fh2EvE7uYBkNFAK0HClUCJ0/wQHGLKdt2XtRHLmnEFi+nxdi3scu2CeI
1+Jd2rlKcAyodA6ITGTX3PWl7Vu7dfvtSrzJfb7dRHr8OmfTvi9cpyh6HSaG3d3lBaHCPfCwvl/Z
vh7ELpmwK7wmExff2WmwrzPD/4oG1fdZOzjXno5hr0mtvFRFwYIj7ei7Rojlgo8SrWdelZA+/44t
52Vj5ON7a3NJ1jqNjexZiDEIlBNMF7YK5DbSJ1M0Q0jRwN/OCRcnyYAi3PX6koXbANGYK+3ooJYJ
1kzitVeHGiZom8/SazDEVH7TcLBx87uQZR0PJ4T/+tH5Sp21AcDuefC5WRaj6hwt6E2kwYyEbjZ4
TsWi+H3gj/4k4J0lFBFvp1J9MSEZSSzZeFK8J57j2qjGIXsJC5/QofPCMv2GocsPSDNzU5gZ/31z
M17e3F3EQx2YBIaSOXuMq5vi64a7kw96jt9xAN439dVuXQy5egCGktZCBA4hqI90PihIZsYQAwGv
L2IetHA4BRJjBYdTp1gtjbkgRvTxM3alHxd9dmJ22B9erKRzvdsZTSsI4SgNyD2Krr3qvLl9AXKy
mZtUzp6l08qOhQBgzZA4HnqHJ2PqZrOyXbbpWzvv7Vz2ByR66k+ts2j62vTc8qKFdsBVtXJDI5Xs
sb0XM1OcPuDXcr6kh2g7oFqFimH2VJ3kxJdTjLiUP9M8ZYTMzkdyhA8fvWOnRA2kpIFUqw2w9pzG
uFjpgHGyKO14BxezqBddM9RItUi2jo+zUjaXonMojYoxCWfFTuv7rG/buU/8xwq0E/gfz1WDdlFv
GS5elsF4qovVnIvol/dvkXe+7rbln3Oi4Uigw4iPwU6Ha5pBB79VmnyQaqfbWJjrm05J9NvRgVmn
ksuC+fvTUZ4JZrOp6cuq+ENy60/GN4IRrQ2fv9XwNJPOu9IThE71NUBRbQmhMgvoN4r9o0B9X4QB
ViUkzuXZr7hSE/uJYPpMWFSTwHNfCDTlNbFEwc2pSG3KLXlrfRJpNajeD0myujQUNmDp0qRExtGO
cSZ4OnJjebhf1y4QGGm6JbIl85G+NUDsAHa9H4XnZAFM0924T8PERSM+mDg06pIXN+bT9CJh4cqf
y/d0GbURaH2KLL0dGLLRCIx1DMCKOLNggqIo+2iJblonaPVdfj4/US0LUfLspJ/WVvqiF4h1jjEK
FkWptWUHssFooMm/Qui+MI1pSx3x+02TrlAfpOH3HyB0rDzkwQjtp/GSoL+LpW1YHT76mY/sdxsk
FV55T/QQPyTVS8ADvFLQRbCZ99D20aAqSHK0mXfKZKsTPWmv3q8QCE3pVhXuuURjpu2VS44NMQmj
jlQIjy3Dqu9tYolt8voY2DWI8ZQbzuJMAFt8+O4u4mYJNJJ1vQ3FHpJwBLKyxVOT/yJlq0ieQK6n
SQ7C66qpysDX4My27PC3jI5agD8bZd20wVEkGeURkRgnk2dCaX/vEFJwqG0tjDVEClUgo7knM7WL
3WFBbCNmYJcI8zquVVGmZsDbvqQgLHXmnDx4fD2HX6i7Zj8eUWMm7r5h+ArTZOiP8S3D9RK0w0R6
eHuw5X2l52fbFkIkW4tNjaXFNUkul8ElnzXBIXkUW9D8TANymoq5C3PJR9UziRQ5X+YEi/bGNpun
PDtqf2kZmiGkvEvJHzbmMuQk7UDczOe/bcGliLiDY7afxcAYiCU5vbM4OUGoyohqbA2PjswfOYQt
2ro+7sYSlBKhD0naE8qY0LN98IBnIs+cMY2JIZODpwP/jAbU4Sj9cKM/jgzRgC0lsQ16IjRBNG+R
kxJlc8jeAnTkb7e5FkAiPmglxhCrxDl8NLfBolv2K5RxqctWwj9jHWHhitIZBjqi922ELJCEex1l
Vk/FXOvQ7jlOtf28tesBuImnS3L7PqqYaEu+SRGmPexwyJK823OilmDI1996kqkIi1e3lkd6tBdZ
cA1LWsAdN8+STrg7ZZbPPX6ms/VO0KwAURffojoFaB2qCujg+FUqJJMAKl7k8mWC2ph5PDf8eSBf
L+w7p7loHthPQSPOoVWNdWZtZfixoQPexmBbFYil8ipioQXifCqUKzMXLAhM/MF8SxdXhWz53RnO
sxFHiDbPU4pt2TuoPzJnGRof+8BcNC56cdm7iBHj6h5Op16c7KlBfx1qJlxMI/Of2KlYJ4DwkaWt
1C9nguY0ZjYaKvfjBrtY6GOO19aYKXaHTvL4D5Iqs46jjLdM91VHcbeReOKxC6Y8zS92pCN48Rm+
NoV0QSTI4qC20RKhW78H0LFUmt+/pqWvcRzSFzD4nrgqtK4msw7BOVyykN92ib8b8474DHeGeJaf
89iFYnOR2BeBgQm4+ugmWl2dcKzIuCg0I7hvDH7HkNhhDkP1LciBf11z9n8fmu+w5bX669PMTq06
EPdjMyb+UgS7k2OcOkfTobLDATDefqB4fYGBpBtzVWxW0gaUDI9+B2thvFxN7pCVjROpmXzvxRPO
y3aeKnEykhffY/iphW4xOgnqI1h3Nedqyd5giMkJeBKRKbigS0nRaqB+FWU64aVVAoeZf5ZlXG42
RItk9Q8Z679wmGifJPqgwdoRuvshNG2GKkyrkyPFtwFiueN/6A330ePXfV0x4HMIr7GWnHKFiwix
yN+qMtG5tFMgBHZdrSD+d9ylVbAZ/aDk1e8VcFApXqgnEIrIS6yruQQHRKH/PUGqWRES6aV6Q9rz
lJyDGL9SPRFt7Odyk8LnWUaHq5y9MLT4wqLdnNbLF5MAku5FWfyKsz8J1vxTFBtz8lRoaEl6P2c7
OQbKEhIFiycueAQou2cEvDpmLZ4DJFqR92JDe8PQDXjto1Wij1kc2/sJyUKFWKZLoHier5pgGy8p
C3woFTpLrAsciqL3Ls9IBZkD5EizHQ03pMwIgp/ZTIzLsUFTOcU/Miiu3xMuEGe3RHyy27RrecYr
Np0/hZxAKwweLWRuPHsRlZ9Vc5EAHgBZIu/XPP1gUvGw/CvW2FRP3+ef/dNmiskqUkF/KbMGgFw6
NqNzdpEdlKbjW7DPF/J8X0l2/y5QuuU7lNK8ndnkhVVUbQrqMafqEILdS/k9wRGoSqEYWwDYRbh1
0oRpzTzb0xkt2CuSUx0pmc5jgewMnENb3w1RvR3qKF51VffeH9WXktdoasaxkHRKAUtAZPcQHrED
eP6xv86+awn5wI5mtajTL2SaU2sgegbPfcVjov6304O87mG294N5P9IxrZ3gAONkowdS+ISfExWZ
vHwMvUmgpksL+OWuR1IMgdNcrhXF7L03y1T8cuR/tpbmZ2e+O8qND3Se/o1an/pq1kGOyj1hKgEp
2TTHpCsmMjheCsDez/esHq6RCVllIvRftyX+4iJ4/Jzb7Ti/eks41k3Ri4fYOlnLC7AhE11f5j8L
kwPdo/jm4UlJ5fNvtIu3UaeGd9I25K7/6hPJ5AbkuIPCsN1zBh6MNIUChA3HQXeBtji8ibG54Y4I
oqoPTcSER4b66mQt7i58/5KD7Za5VZIRD3/Trq+oK2bCZTwglLcHIpEvByxO9r8mPoxu20f0wzuS
4vrrtXyczt+WV0/NKT5U3GgVIY0v66qsYN6UDJRrVnWrUCLTll/R3x71LXmN4vpD76h6wF3GCDJh
DKZ+0cbAItLyGpw1D0ZkN1jMCEo4cTKBlYZjOYdCBrymWogx1r798p9/nl9ZOs2WS1Oq5tICUGqt
u+sNBXKayKsSgmmBkgcyrQ+U/Pi5K3azCuqLHezsu/XNRkgSXhZd4/GGmQoxxeh7VftR71yYI75c
c3CJj1zralNF41QJJ4gVp9meMvSnSBTtC1mrP/wjF3k7vx/UmMbivXDWUb3SlNZLVfoFuMtvCKbu
g9hNy4X5m3RtL1MFpWyaBFszJ0FctwJ/6ZyxvvDoA9rR+8bgcnovQ+wIMzsBZ0DHPS1aORXjjbE7
JIl2v0e9QYYYUOpi8AhhaPfq+0aQ2TE0elHTQii6Rh2pEcoFX7Uj6fbgRCyQ3oxXON2th81uZPBY
NxBQlCJCxbmZdheL/9C7Kw2yky5zmUR4fjTknyWTM94sSTL/oKkAoQYzumkZxAOehIL2eZWpJM9B
qdhBOBv20E8EzGWDAFrTTXjbeFVG2w0opXvdkkc+jEE3iFpm82zR7ZXMhlFkYRwWLpj7GMkGGkTY
6q/UyQNlLch0V5KFZGWkjTkICt4ce8uphMXgWtVhU/5EkI0XBIcoBXI+wPa3VscqjBDAJ+rQx/DH
gQD6hMst69at+b2W5wP+kkBBeMHBdVFNyxY+lt2CvFsdqKFYx6CbYwhCmj+C4OZHsXRaytQuteLz
x6Xs+fftHnnmduM9JvLPrOzAgA8Yjd8DZB0YyzPe52CVYyMW1tO+N0Sa3/hpc2o/HXCMnSnBBM8l
5dCr6oQ38wybXFUbLQcSijjaapZF4Jxjy1tEE3GAjQMT5DdjAmNwHQMAl7H2LE8IUlFQtXuHZsT3
5FDTWEeVnLmxnif9sH3K1qNW6I03/x/+UJi13FhEXe9j1dMeYGORSoe5vD4eVH8mxjBCrm71SZ0L
RbcJKOGrz/GVyLkq0axz3NpdjXLs0aK/nb19Z+VvGkuzJmwDQhQRPgYrhRU+tvBJC2pF5Zpda4Zf
ZDtPIiEK93DxLU+rsBwbJ7lIIgOZSs80bRh/vIxYMa4W0SBPCXLqKkLHodFIqF46icToiqq9zaVt
vaJfDra7t3DCyIdw7Som9mjIayQS1p+DWJRvDm8HknfImjjustpe1dAzhEZkPL3/anENMDHsGe1f
8d3mjFFgDx6p8Qz+ONG+jfRSm4tSnDH1eoWVTBLEF2mnjXxUZ/7Tb40ljkNE+bBqNvqTnTPGLud8
m7mrnpSejh31dkxgdz7JIfwCUqw35OnxoIaPsIkWaT2xXl2uqX52H7qzj+mIdcVHqhoo8/Hmkysm
tyvE3aBvOu8gJ7xzk3XTz8PeTaningrNjsL8GcfUdG4HpFhXR0X4ZkklCbHzpb922LEzeKncyK+7
zxISiaXHbxK15oady8tMyfT6NF40ibyQFQaWWOSyRA6cQjpkoB2KhH1GhqORwAOWchaMDkF95unL
XBIOi13NurRGn94x/JeD+iMV2jMabQumzCMgffT6Ki9LHJnTKn5X2JInTwKKEFb7o9TTx2ON9mIW
Gn7bpPQvC2Ggz/iRyZ2QZ3D5qjMTg0PyEx9el4BxMFNBYANSZazJe8g+R/Kb+648hJ3akPbsrwfT
cIGSmFgBNF+eQ6k9V9y9kESAE/wNMC9H+WtbxGf2FodiAbP0IzvGroMJNSI1KPABbdQk3gfRWczl
8iriuww8/+d54STes51/LWv197iQ5J5CV0SkD1YVF+wxKUTLZfmVicabnbR6WUl8jVhLVqsBbUeN
dHu52VKfa826Vo9j0WaF8jCD3onAtYGQ4e2hidvwT/W5ys6P4l/mmnmagq5h+KmIjF3IySbbwqfN
vEhdwGvLBRj5A1wvHMiEkhBFEAQGASzKNgvfaEWgMfCxEKE2TUprm6zOGBfi0dEbXJru8Rsmffln
qL6U7bNc9fDIkbzBQjMz0JBHwNG6lshhS88nkiDf2Yu6kQLYboU5XKx4faMcWX2zhhzq84755Cox
3pgoPdMd5+uGalrpCd2k2rHcQvyOCnvD8u/ibrD4+cjQd5hcG1I3CDfOuRFSJfb9+ZW+hirhv2bB
GmSH1+KJaip/7XGgu+YF+ZwhSkiLhvNKQ7Kvnu75ra33WyYuysrjxxkgpZWfPXIkpzKOV77m1MbY
XyGWAnSNSYcBE6j89p7foAJfLreMYSBnFq51oKCpwC2ds96f0k1geqeJ5FHTBWQutRcBHNqJPNT7
tuYqBOvQJP82DtNqsZbLPw588AOnLSNYUgbQ/LTnpaqHtUS/1nbZfd43CKtymir8Xkh8X9PT5Q7p
DAZLFVi/L7YA8tVcCoWN4QkjJAGoVmDPsPSSe2Fx7NEX4a2EO46bAOpKOw8FPh8j29V4TjYiHIpB
JNghcFCmP6XlFuvx3tJy2BWelMY78sYHykhcqcv1KXm9q8xNNkRkNCRPAlADAaTRLyBAD4lr/fQi
j76BWyas0DjVv3ep6q+t1pqwElMwXV8C06OqmEW6cb+045LesfU8WAVVYPCtYx7Q7RSILSqahyi9
85lfdxSn3wlqTwisJ+Yz1QxToPH1B5oSYERUCD4YWqucCzKiwvsBh745xm7mr8wQUTv+jE/E8uH3
Osf8wWO6q2jgmHYC82gOAVcS63TguppRYWUioIwi2Ef6Ead/1X0KRAsbpe4rR4A2XRqXeMw9KDSF
EZmpIukKFQYCjxuIdg7E28Gz+BeTMkNvlCgLyg+qB8pB1gRhz1NqofMmom8HHMq+ewb3WhO45KPl
gyT9PlVhulWbxzzASwiXQY0iz2Btu7pc+9XLs7fPtP/AlFMamlz9PIOGw9M+tq7huKgUxYgMWf5i
bwmYxDYdr7wzMo4LcIEw6qMHBx6tnihzwjCIMC9kVPEGhjBLTmCqIw4X89U3nGyZFtAurXb/e7XS
HaDED5188CUcEjW/Xg+gStu9YVaVPtd7HTrCmcNQIby8qIpSJzVrlLKCRZffw3oyksZwWH1x2Ey5
pPYvUZSILLYCKIeOpy3ObjlTRuQYH4S8ftUDKNi0KcFJwid00/7MT51bNty4gprKW0sA+f8ClELM
Gga5vrkxxOPdPwDkvAV7bqOS7SJ3lBMs/3K47Am5vUEdu7bHfw11uRlbsWj0TDfyHUYvzQYrWJ23
THeAcaw9DJ5WYzr+1BnAA0WeZYH1R5Z+yGQecJn3aU3ljrYLMVYE+nisCcSbihe7D31KRYMlQqO8
fvvwRtyQuofVDyebA6jvipUaXVrdkDNvyV2WYp7d1OEe6Kd8SQhhJ19oMPZqYyvzLVtwX3Ka0bLJ
OdqK7L643LHqAFFLj/LDLwMtHFhJMR7ztlfaSiD1AnnqnLi1Kf7Z76gfoLWgYkLjyqTFZ9fe0Ytr
fWXl66SLT0Bf1c+xObMW0qeQPz4uZRKM3RzwKuTlr6s4eKttNt6Oh0LogtGySn+5+WYBqk2jCIVH
ubarazzSa0uZMUNkD5SAN4y1mzSKNd5L7zwqAHRU3iPT57Wtam75dX/JQeG/Z1X6aelSkaqa2S2U
n63zSSj+xl8/AgrlHuOYu2RcDkZNd9d3fbXzBy2XSpWA1iBqyuooKaBZDz9QVG8oDOSlbzFA++9+
8gJ/60xaMpVyY3sxbpPsjhZAtNxnbepX8cnw69A+0lTqRudCB1K2skGOKM2kHO+0yOgOWKsYsaiy
WpKXsyQ/q4XelfcgmTCq2ZcIx44u8HCKYA5656w/HEB8tq1feyIasALRprJCK99R2ncgav+p/KZk
TXIWL9n31WRplfXTNu372kdtFWQASVBAhSlwDW5pigBHqWt5JlBJ36tCeXZZeMzCraMa8qPy8nua
EgBJAG47PhrXmRfAfyWPMr2DyW1x0t9TmeZ5FUeAiZnqfBWooAdzPjOcFoi5B5xWlPXtFWf0dmJJ
U5umVwGKtfJan5PM7Q4oABUTsmFgh5ZGaKiejACn8nNHAJKgnsY7gTLC3ROhcxjMkYPYjgrGxXd3
B6e0e6RwvLqw3zaz15OmxYt6u1GUUMnvMToypU6JcPRCb/8JyZ7wZwmKRh319KVes1IBMrOugrCe
yM71Q9FGlNI12H0tfFacN9HpIM5yd5d93jlr4ICzxuG0zXEj470YKYDrK2Y1WapNi6Xnvosbjo3f
hTSaKLgThs2PNssxki2GsLkTKi/6KDGEOPco/zM9fY1nSAvxV0JGd2zN0Ji4YM2zuSjPdurFn0S1
8jrlbpRxi1iNM3x9FvATpivqdSz/MwVGHPcD36VSbRj9p5mYo4kJZV1G8OXGk14iL1k24cEECPIZ
s5OOIYl63iSlsjEDgMH1Q+PV7eF4NM7fbY4UtlVpetpoVRNCtv+yb6j11E8CCCVLA1TTBJHDNZSq
2IFeAHJmIQaDdA9NlLcAweEVu1NcKOq+m+MKlJmO6wcAxdJ0f63bBMh/4hTQgNK+fWuZ6yH/YFan
F6A1fUKRu4oII+/cYYa9ciejx6oI/A44FotFit9E5Pz/mz0WlZKCgF24p9G4AKH4a74oFuWTk36V
o3IXgHihxDMcflhB40Dwb1AqP8iOD4PJr+UUiC/cySOQ9fjTpy63Sv4NGeWnAC9Q01x+nteKmarz
I9lqEMyYQ81JjzN1MsvBb5cLmLRWjvZRnV++TYePUXp7pTImJniYR7ht73M29RdqC6h+2AbuZmfZ
4JNnVf6RkJbkQXTSrdDt2Hpq84VzQGJH36TsYsUuwbipwO/HvjCYOlPaoVanyS6eTtaj7gcSrMSl
QXimlS7Ral1WRFS8yZgLkVdk0r0MBlPywAHXTNlHJwykhLlHk5N5cBlhPrttXSy+kGkqxGaoYC4Z
csLVbUSfpUbgGhdbuAm9juKTuM/dFXS+oIrOeVZktBNVDevUg2gX2BTXaK35Ba5ppYdVA5lskmbf
oHGIqJYXN6Oh0n8biVRgwH4f0wGiqXS+4O4p9SouArXSyirxJBltlrll5wNCUuKVKPhdiWKBJ7HY
HmYuYmtY+zMgNIQYv2q4QiVFxB9M12sN1WU81bf76OdzYl8BOKH50l41Gcc8t851IS9x8sXQ0YkX
cxhiBd8hzIdIucFRN+b1lLu9dh6Zt5Yy9mE88Bj9f1mxbY7HT1sp9+UDJU8N72y1B42/n+/F7JX9
tSyS+5u5Fxcyvyh7+HpIRO1AZzW7mga/dSAwZnJlsZmFu003Us8DHCxbVE0IyNeqYEz7tMq70+Fh
vnk8VmYlFd5x0PY+Dr+Mg+tcW8xlkdNJqLfl46WBJOLspKKO5ZhY9a3gHCu1Am2oFPYcsH1bs//z
YDda4aWXSx8K1SFGTqKXyVEFKNSDtzwGBo66ds4ismgFQs+7PD5bkV0FF7M6qJgcfEbLyYj/h/tV
Wsu1rX2q9xuhgL1qkJ+mbUS6XJYdfRMJqrKBc7d76Oebty5ekvTYEG6Kbti7P/ovjSUn3YjsMxKb
2G4UiVHzV2IhxsdGqjrK7qSkYS5WI48ydv0fk0Lp3e7SIGB27kEW7+S+3qwuPdt4SmjoKSXuuY6N
zbWbfCwaGlKq9dYMR0fdgyuDSQOKbCVjvSnvVYDYhAwP9jYv6XJ3P0bgUknvukFDcVwgSeouL6S1
G9g9QkEXlZnhMbHoynfqqUq6pro9thazfPRxBmUEs+ka9wD6D/5Loh6TfbWNmIi+YGFG/2WZqYc6
paFZgd0Jx8bHhGsg6/ikoZ2lBZpjQx4ImXE4iKMffFknsgrCex8CQG1FSe8Lj87nXmWjjUtk6Rsa
27AlCLwHkO/YXA25V/C3BW83FB+BjmImp+FB3BPwKG51cDGlkSOU1xRKwaKlUfb/1NrnV0pMirSI
y9JpJ1MVNBCymZz1Z/lzWBzgEJR8aLuEpI4erM1b1WUhv9Nwlx+hue2EdLycGoV348WAYtfpOSy2
pTWYozabQ//8u0apcASg1oXmUFnnktY9n3KQ4OoJOnstARswfdTuU+9KuCsFi3n9l+BKJ9E44kvc
TqgGHPOYn1xaPeGfsSW0/S7+w8qWH5WaWUCt6x9OSqvMMUNQNorQA3ajWq96Ey//pdE7ru17Qb4W
5MxtyYFfP57u6iAQpj4PHCdsn81KedgI/gIuT3JYhwYWZL2+jnx8mFWxKwexlB335/5QVfeSFYHa
UtvqULDHWZGXJvsYifnvzOo0pXiv+qJiHkOjVqLb7qFtbRgqy/WOuJnUTOcjMAK0NcLteG6MLBHU
6JcGUh8YvG5e0wYqV2cXOy5ArZmbkHrDKJSMAQgjTkDzdA0S/kF67RYkjkYc5zdH/dxIzLsek1oW
DrpIMqhcN7ZjeaO1YKIki2MAAPNvc+ra1IBmZ15gGqbIZfG5fM2mOkYT5FjDu1CZDAdsj7Xy6uH0
1OlB8zcQLcWehN6kb0LeWpJMKV+VNZS5Fm9lhmBG8aAvbDwYshqQsqc0h++QwvTQnnLZPd8W3G7P
6r4OljZ7wcPFVD3+00JDSQhznmM41+tngUjZpvA8FDbWCn8JucmIRbggxN7FHjAlQT7LKypKLUbv
Ae+lKH9BFEnBIeSGfoyRYPwjsAd0vu4TmC7C6W+8SqSVHlTALiTqOE4+Tvc2q8mkdSSoza+EON0l
AFd60gezDwmpzGmv5k5VnW8TkNGuyF8RNnXRLCBIy9xlAtZ9Uun6zP2ID6e5IM+r/n+XJi4ZyA1e
hM7T/fcaQzTIQpHBqdRfTYD3nVmDNTokt+YT1Sy8O3XTLkJbZd2N5ZxvSx6thxUSkTA1FNPm5LKU
Bi3bWcJjkKvAh3hz5dXSyUTD3mZbAiAjTIuSXm/jg1h3K0dUzdwpVMys31YybQA87UxMxDi2Pj7Z
LFL7Sb2wMGXh9sTxspEUnCnRHdn94pzbfJpHmJWZs+raUFXhObQ0s9O0zUKIrUni6gj2fxWQOPkL
sv1MRzBULiOlY/G/xjKRTs2T3mmTP5E1m7QFEtM6mq5gbaRAAq9yw4uc/zJmZMNgpvG3CCOw19hZ
jgRvugU/UmqkhlATVfgkpjZ0WLhIsa7f5i9T3ixLNPh7mWcwbeoY/bnWW+FmSs2EuoHafJB3uHSw
EffsmEHMkWwkT1gRGC3w4XaQ0UUhajcOZZH1wh+MSi8tHXghyrv+JGszHuNvSsO0z7HB3qIdoh+m
2NyVitgydr87xhmpfSS5mXLcpy67ZjByMquHrMLqk2/RbhyMJjwBNRpgmz0NCK+CSiM1Qcdv6uBV
+ldnNlR8uc7llfLGT1BLkhBh+1SrbQyYNe2DUWCVrin1GJsmRM77A4VT6ohFqu8b0wVv+cPmwVQe
QnBe4pBX1cwp4T7LdUnJE13KmU8n+t6wHv1CR/t1rHdvOtgFH6Mzv7EUiSr+v2QSytUrOkOj7tQ4
m+ZSAB26ZMqdQlIxkrfAg9xygdP298osU2E0BK1sF+MUEG+16beEkTxae7wOpNIePcoGehphD5kL
mxCvb9ls22Ikjes9Z6wD2A0G6EXnAV6xq2OaSCRmbu/Ru8yDYYXqdPs+h4614m6i3IHFmPXOW+DR
G6bTlsMFC2FnFDQo7GzRpVTv/kzUMuW4A5tDdbOTK7Fg/K1cQ/LcjQBZkdULH4V/HrXspN8zatRB
Q8vn2Wegtw8AXMiWdkghqw//qQeRmy+mqm7oUdX+fdbXet6pz5WynTf+fGFW0wk3os94IbtFcfSG
NBEJ0xM94Us63vYe42KhvTQICpVHPMwFwYq8+i23zFfS3daSjyqU760jVVmddFWskeY27ny015dy
z1kWGwqRQAnAeRBDF2UUBSIst2ueafkO86jd+nDOafsjTw8BXFn28ZhNEhMucFao3WXOHM6F5iRl
AYoW5X1JK7jihOyLg4Tm7Fb/7N0yNBRG+K1ysQb9EHeQofWW2zFpi2G51y9E1WcNS/dHTchxMUIC
9Muh6QWjpohV4RUOLVYbu29j0zWEWNqYtL235KMIgNCQ4JfBOI58u0kC5XN+6ty/fCS75JW6T0Zg
WgeBUBMOgD+xJPl3FjyfMA6IQGQvF0sfwcVtPFA9FKDjJYBi1CTu+VQqycRsqn2zgAITGBsNk7Xc
27IuAFFjvppVttm+cZof9+vfDDEcHDbSo8/C2IzPJROE2ANivcq8vrhqhrKCT5xCe+fZ0FmQxLHJ
m87CkbMouTsHykl7+VNMjd+AiwZS1fQwtjhS84scqpco2FWTw1nxyqo63f1bOcXv61v5fmpJcnc+
JJp110n994DCSfouFih90x+/EM1tvMMOKNu3dzP3rwG3eVnkLbADcwLmTgGwXACp3m19YVZ4cD5B
fdgNAWIywjSgC6Dk5seY3P25jCxfUJkpoCIqiW0kh2Ho0FzFdvFe6R9jT1ARL+q02T3EVr6tHEYE
aAFFS4nv2zdDb18pKPVQiTRdhKlQOEWAlZsGh9HhaGlskN9VdWn9+Hr9GjiOYZ5bYF8jhtWeA9ca
MDnxYggp1+GBZdaCRSqs37O/+9l1RMg4mznHRASGZgjhLVDLffJwWX6fTle9MoE6PKd08lqf1n+3
RkO9WkFDrbmJhXBoptnxy6GWJVxW4szvnr+OaZQgcZO8XkzR6CeRPR9VmIUEUGJBcQ6FwTbFHZa7
uV1nf2/rj1qIQVUODq/3EeoHlCZSFPLpRrarqzrwtAhNh4qxYqNvsSJETZ8SSmZI7O1iHNshQapS
oRFyVKqufTZOiLs3EN7VVry42E3bPRvtyYmiN7vHihemqpe83PdaAJroClEiQmVtWaxth37Ejjca
MDaur+mEMwFOauzbh2Y/QM4L8pmZpD41fL7v89PAIoqpD2xPvWpJ/2XN2OPNmRtl0dtEv5WdLSxw
PeZseuVjwXcwsgicyp9jkcx8rSxZITCk0kyA6gVPMVSNQ4wObZJhjK2Kp/p8GG4loa30I1gvDoQ5
eZUfnd0C1COOBkkbRGVpSKLBOw+Nnj19Yw9QcYRaGaO1F3/RKePgj2Pb3iYRE9BS1ZWih8rnPIT7
DYlHPRVBC+SpsLL18a+aTpDHzkBAhaKqgToK6lVk3Zr9V+v7Wm/4W8Zi4Q0lzgK+Da2KU9orXaxw
iGhSqdNzqNzyRSX4D0AJbkYxoUS5NaLeG1FRJBiaynxpHHpkCydeATBPhDCaS9A7TbqUBy9pEh8+
nJ0ToLJBkWALGoQLEdNHCHcLiIxqUTpknxj1+U19OXq3ZinHNwHkqq8IbFDXNKDxSOgrwHPRJZa9
/vPnt0tX0m37iDs4gcfh1+5IPJGs3YLVT1FsVCTspZsmx3FpbidZAJDh1MDCIRJlzZmXtgTyWvsP
GcHncRBAZdRAQ30g+psX+n7ZZ2E6j31cSKa0VUZoEfUpLfrj2/W3eLYK/6HXijmMWWnTJLnnKGPV
9BXc3fqWdpzMfiaTcTN+XsLRGnHnz5p2Ppnugn5aisy+Sa4oMqNuzHD49Q2CgItNlrTyyXMrf2Ak
f7Hjm3vdSnlOM0OH44nYseiUHSsWj5xe7hufWTcsF3rQ4RgSN+Kget7L6YNJfUwG14mxDRIlrjWJ
vL/a6vK0WAvrY1OFEgglZkL5nurtuXhmefKoQYv7Dk6tBGu8hsVuUiQ14kq9cdr9nA5YPR50Q04N
B03yOcyyiotm9DMSmOJaEctWxKTHk3bMBHCnhYYvMiNQEt80qVla+3GR38hn7TGzQmTsPPHh0wSp
BqyF1bQqEEYKAnyHxXRhvbiQpUiX5XMc6JcWLFBc9xZrVqGM/qVUim3t8W3uElLTYqjDcl/PWEy/
NxdqtLCYgqdUJ0YbwKPRLFgH2VVF7HrjM5Fm2FtjugUbGpabBzOxS+PrJ1P9taEG5LE2GQghGo1E
FlTePijzcFBv/f3xNqNN/+QXJzY1z8VX7CVXMt89ahdXPS2Twg23OygdeR0511KHWg6WUmp2WelN
yWA0u9xaDWv03bDgSDD/g5TyquUELGD8R+JK32n8teqaofv5KrikvA53FwqJFpGVfEZg73rNlUsB
nlmgb2QYnqrRCSRs5shR1sVa9tIrDWZZ2gZniEAJvCrXPr3VqDPkus0QmAGtnCclshV1AszzYdh8
Y2xmhyilzqmQ7niJ6LYZ5iSHtlA4MB/hnb+nLBPzkaMPFwQLv+AiT4ydISwQFJtK9W7kr/MbmPKJ
5ePiRg0vBwivUdQptsdZMgbEJE1Pyg41WklKM/bbFKGdOYuEt5mQdbnxSz0wrb/9hnGrEdKJrpVR
SB9G6UUTG9Nr16dyq9Z/+3tsS+217XulkzNzMXaBIY0yEcDcoWySt7qZCRVoHpPEslQE4OxUOyVh
yK28I5Mc3wXw6rguFK9/j76ByYAcN5QwOcaT06T11pC/jnyeepXDxGzBBFkdrkGX+pFcX07PmNeF
Hp9/pJRXbSL68t1xeAmDR7UFOSb3M6dlQBCCLmZCnXkzLxfb+ZjNuxs7Wo48+e4FkzTEoqeHGvz1
vB4NJt1q+qUojYg5P71YklQHlXJGV/YgXdwcxEOFLqfgAg/Yx9t/AQTMXCBL5+gUun6eXmkZI2XY
YqvtzG/OGoVRk1k6lUz6BRgK+2Upqwa5P3CNyWJnc2i88SpGiCVbL9kVxwV9dteJOrfGyokepmVM
l4/ak5rVhQgSdvZofR+yNPPzpX/mu3QXKuw9Dnr/LSil4unRMoQRLPcaE0OJvAR3/BAwupUhW2zP
EZfAwmHR/fGD4JD7lgVyMEJv4hboqOy0jkweXZ+TTGTXlB78MxhVsjL6yYp3cS6Xa+7Gz6jDDj7L
+2WmNsRBwUev7ztG4TZFHpsqFOiRaBQb2kFUn55HJqYv71QQTm4GE5yg9bLpoJ5EgIYNvebZrT0P
ygc0ROmfxnrouaV19yQWdCfYdZEgfia/zYvwngfjH8ZSEDiAESeUCRZCIE6ckbzB0OthR4gXPfzc
TFOO6GeNHor3gFj1KhfEALpRA8fWSHY1yrHGQpENjXWIU9tnjwzLbkRHMN+sO0kPool9SGxPV/8A
B8shLUYT7NYAZXajXhqyn2zlyDztI4ENKvDyKBLnf4DHdMbYMQUoO8sEmtzpE5SldXaQIRSEdAm1
7uW6dJHk3YTFNjYKSe9mvThIxiIBB1mYXOEFQozUpG0eZYQGuO1WbR22zdsL+rwsR3+mh1hZP97P
yAvaMOGukh4eNxx9xDggSlOMGDvXAJkDZ48pZjYyoR5FF4KwjKDN0D6f/umkdo1PKtO1a/7OXYst
roYfr7m1UbhautUSPeZS0m1Bm5YtmSKnn0oGmi9K9orP+g6RE6JvHxARwKtSRi0G8DoTSf4KWHi+
06ybDAzdaMXuKtrohGW18pp8fzk4ISFpSDNaIa4ObVMz0C62YMmcJZ1pDvDrBVkHVD7vk+RMWCF9
tp1O5TXSr7kqyDSRnUHUd2obdcNPjtdw8TkH2ZnUe4hZLJ3o1n8TBtxPs1ioKpMDGQyrwggIREyW
HVk68ljqBVbNmmX2Cmt2XzWiYOKTQcrFXaJxROtPLe4CtLktWWOiv+smu1a47XQKhWWLHj7hIWsG
vZc2M/5zP4sXlzW2MpYVZt1AJ0Nkt586hf8j8W07hpC7sTFr9ZRESTPWr/58vqOljIupaR9QNoHZ
C8v6pBj5dRj0wVCiMzNmrHPmlW7tpNkImfTKRAtoC85haWzGrubqGQnyQmaflei9RvKYDbj/x31t
qOI+aR4U1wsV7qX94YsYmabjD353JXbYKHa8duVq1puOOzGNpTz+1ZmV98/a0r8x5rizn3NDubMx
//0Nsf628iQzBrOuzZldszfWvEilk7yLAFBxzRE0rfCZm1AMeelvesxb2JwxfIOM6GQ6bK8ksfy0
20m+uxETYpYWgkeYHXy2eW0MT7Mzd/XTcBbu4O+M+vZZfXzL1eLpD0nsYiQj7OzNEyqmyWIILUQQ
uhZpsy60wLMGB/fy1T/wkDwUsrYQPlEdyANECv9+cxUA/kCOZ+gKOn+G1ey0gAfFFNJqxgbGFybd
XGEgBhoj8kEk0+m8oRg7cy6LzV97Jrc9vVK5Wg9t6IZKfpAuB2oDn04PCGDkOtxi8rsgsG2zCFos
9iIbqVVFkBZqLpF4mievQ5AMHUcAcStrweb4t2AWwsYLkFHcnLqf0xRyM7JcdZFvcJ5+S4P2JW5z
z7poD8h0IxN/HfTYh7O6BEAhdiMp7TIvG3uJCmqwlxjW13i2eeSE5H7PikoAQvWhSK5aalfCpU7n
pNlWeLJdzXydtfdZlWTrUJqKuWp4saptqbdnGYch6ZIW3QupKPc+VbLwQ3Cxi9slopWBpGpkPZKw
mTpV/yxIXptwGZGO20JuPhoUjLNzGRLkMgZrGvcKim+EVQ3ZdIFZd9k6g5Ewpa3+CNpPwFGVRK/Z
UG3b5FCjSo0YLoOInSotJZTo/9nq68HR3OEZmWitVde/2MyjrJOSjlqlg+NCu3ba9RTWU2jQoQbk
HTLmHvhoIg521Vp71zTYkCtIO836FDWFBs2ywd8sbhCWCzDvdv31t4Cdui3c0uZpAzgv4RwJoetU
2KBLQcDzlyNdZFrhnDXAzxWGbOdNZuz09vvFRs9QNaYtjMfeZs295xJHpmvUSWq1mj6Dg06zv/TM
oclH1YLwjxFHreV9MfiIiHfTkKwLj+7w01Dmw2+0T17iN56zVo9gLbVShENnwagouUu3W4dymU8p
FambKROsD05hufpvbqSiPUI5Rg5WgLi1VbWM41pkkeIRnvm2KePTa+W5tHxL5JbvTsB7bZQHTUpe
mZHqF3Eg4hsd3qxIgiCO+yigq1W+dE9JhK4/jNfk1syTrlDQzlvsuHkLeSOL256m1X47CXFU5w21
0rPWg0hvju/ltRJeRwRq7wS2fwS7AkfDheSV/kuHDohrPYx/IxrSjvpAFDlvc/bjBIPtcrLp0tWc
mg9Vi0Dd1rCy0v9tidNaIaySSzTaygR82kYt4aJ8YBoLYjj9WOCzoy7NkIvSzOrwpQebO8QgT9/K
+S49RMM/gMWWUuxGcvnkX+SbeO6JUglSEg7kejkoZquXdet4VppigeWkGZQu+V6XPusRucXqnu6R
aMPhEtYuCWX3mHTyvFX0+egiX9w18UAczjRCUgoh3C3yg6upmuvEu6toB56nvI4brzMxJO7HymoV
AdPdsuTrM7ROld+4DJ0xZwWqYc+a8JQkrBiia4re7pH06GjPFM6VXsz+wz25/iiv3Iy8mpfR8tvc
7sBsGZua9Qh0/zZs6P8UB9xfoeKu6Z6pUiQIThHkRwVubIGf9qCDsWFxfbNgpvofAr3ahrkcaT1W
XH+9hrXk4WupU8TWawd1KB6ZHNPPb5ft9q1vNSmVYgVXHKRzLC+GMRLRvn4C1EG7rtpAmZWUQMv0
0O5yysy7kp5Y6i0rC8qWALxMUDMBIDcg2cD0ujGU5VblZMUtmA3DlmVCG2QVF+P7o7Nel4b0Tukf
2PEw0bl9Atz0KD3E8D/M0jtYFXcwRyDCLHR2Z+dxoWaWBR18k568SNMGW2jSzgz85yqdIvIS0ajC
kIyLDFozKnr+4NKmmeAZSmN6NkPNDe3N5C8rcI24Fi8YLcSuUbT7J+fqUU6hmimOFDWvgbCRBejf
O08x3r+MhnsdPFHT6PobNeitBIa7Z5S9w+auBjZESwL3xh4bbrSxGctXo/UJoTdkAqJDblpnAJvo
prgJLTc7faBSSvJ+sWX5w0N4cw0HNj5XoVj2ujW7zilY8+PnChd7nszeKNP9D8TW1UbN94VFYh2j
shm5nd91ukIPUxitcXyIqluEcJ6bd57ALbFhtQ96ofEyc09cEp4rA74zkhpeDEq0zMUUKZvvuetx
iIGhYjLR/DNeKNSSnRmUGnmV0p3CsogEaNis1t4Qr5Xvv3T3W7ee7/oP+yVufxN9TdOsFr//qylz
DWx6iQ9yuU3vQmCXAUVN9ttqqqswnCieSENdjDE6CNxVOpbV//XQFX37moN3L1H0OegUuH/NI8Ka
i5MUGBNQbtWNb4jYIs79MVnno5SNcWKxOKz+h9LOvweRFouEOk8cgkLwxUHGT8vboVfwbcvpeokN
ufzjO6JIgGuPNGK5dtIQ2w93U/J+LxW98lcfw9//NIEGww2y60dridqfl7Tq/Kbivk17OurMLFCf
jm2HR4J1DPfqk0uILtXhkTB0HgxP1LlLFcThd08ErXte9J2/1j540TdHxFIh2knC5YU8jmAyMwjH
6xCZn9SgW3yW2wDL0E1L4SMZQATnpZbcnrKzs63Y6RQQhqBE4s/VRDSqMxnFIQhPgGRmyv7NCn8s
Y/hw7xdhGfboD0BA2XJ7sSuuQReMByFk7QdARKUoPneVriZFTrHq+UjukzgrtVMliGRrppx4Tx3I
5Gaqi+3kzHkxsVHMAEzVvrZMbwW8AXrlu3NZwkVAhZtObACStb7j98QfY8aKkq+VK1aZ8PYbbIx4
U/+wh8Cv8kEgtJWEVCWo0+hvw8EHkwYObQvnwqPEO/UYKb0bn5AL6AZxYCuzvvvCkR62GhQwcaQG
KqmUdsGOXftiA6yePYKaQ9NGT8Iy9/Q4srs/yGS2r74warZxYQFoK3cRfUempeiKdNBqanQPOK3h
tWUHiY2ikNRQOsuZSigYxicV20Tlfn6sgwmBOhpB08BV9E47q6AIWCIFJ7EAkPdyscOQxe0Xzym9
tqbBARQou8Pp/0T/ihimj0N7B3ilhmTktF5jLMVsco8fyAxV8+Vo6GIz238+mz/sTau99myGE+jw
hxzBG3j8dCBppIGobVTowJcDyCWlmHc5gOIh9DoGOVL2V7WaBt2EN5fTapW7h2vKMIGoCAKct72j
7l1orYibyXzmGoIhl5RvNXYw08B7gYjauClmAS8LI4BQ3pCAh6M98ZIa3N4qJ/9W9l1w1QWFA4Yl
Zwnh/RAnHcwe/Nvsqha7bPIQCSFLGCOAfyUaf4pQ299EzFEpCCK/om9C/fSA/jF8QL6hTgI7ovSD
ttJsQoDPdp+2b42+WfPMnfpRGCbNZsFG7bLF1O7NC9jZr2z9SZJ5KeoCAV5xVAHmlbZ3SrSdI/WH
JtekxYvbdJZwURZKKKDdebyN3e51gimLpiui4ez2wZLm19kx9GjadlV4v+Kb2qyxVoZSpj/TXBk5
sNz/kiJ3Bbid3PQI+9M3VmeAPQ/rB+6sE3cMrLL5+KnBh2xxLepPWeZGUGxsxCwcOuFjTWTjcZUB
aXISso+Ivvd+C5cefcJ+2yf/cpI5vyOBvSulNXvJ9ubi03yPwomOErS+A0IG/X5L3s4axnVh8hcM
K5pZ96qHPH7lLHlQaD+gWGFLaOYq3DOwzlNlF7YblFenNbdmMaCVBba0xKIhZUp7XXy0kofL5VSN
W5ekifvbwGTVX/o/GUv61j7dzPIlhpi328xrlsN3QVQG+oy3cpr+7sGCdLxjhyNhNZgH2ZdW6Rs6
P6kyXfuuc2lAVZcvb2s10wBdRcKd64ZZ8QfeoaauGlJaFItCW6abKuOSU/lkdNS5ZORf6F/MIwIC
mHIKpr5BPiEEvjhMf8cgINq4NNHi//uHkrQNl5oZ5ITEcNPxJUF+W7e1IT63etqG8LYLo1IbLn6t
970HAxeJDFdfzi074+rvvLe6bYrJK3mYvDRwSSeGo9x/etYdcB/rLN31DT478t7Ph4uF6byXYsN4
RU8Qc08Qdqv7RproePrqIrO8K3riigEwkxA6iEyK7qG8z6XtY9eouISN0I0ZPGza/uykkAPUQ6gs
AkKt7MzI/72+9ztI/ws7JudZ8HAA6wMo08IhwQQ36pOTZ3q1a/qysUhd94Okj4NUU0WsxRs43i1e
xUSGzRTqTg27JHOJbjmRT+AhJuDeCjpxXMcAQdLPpxb5hgwF59RUeJ7eTHBfgRXDDff88kz7T4V7
LYnnL1aey9hES821TEAR0W2XAaChMd6pmoopb5kFddNC4a3cZTNFkYIIrP2Eh2PK1AYteVEgAu+6
VI0urjx0Gb4Kdmv4TA+Ti/SwdnhibMJm+C+Mh9kV0OHmyzpo0aJ5zOmRq3W4OG051O3cyWe40hkN
3z16z0sbxhHsaSYQ1+TtFeDQuodXCRjkHodSK5+PMxiktaSkoKm4v5go/iYPSBmpx+D6OVVpBLuD
qP6fI3OHGqpAbcmH/R34vVbwE9nWlccd0WOP50EgZqCf0e3kBBGuvQlTnvTGjPx+/DOWytTbdNl5
HXf7on9QZHgrpTz+7z6osTQMoaA0sZT3cTERRDZpqTaAJ0A9/FNk0BcygWni8M/CtbnWtQiDCUwZ
8bvzrYcBsPD2YEBuaG9RUyI8oqbKslgNIHSf0xLu3RWhqdK941FZXu3UkrLD0dVWbGXZgJz06/cH
9DExlR5HNrxATFi7MVmKhfjrvcleUO5lkeef0EQDFVdemaCDzt2bHs6NDY4ORnTcR+vYPunOv2ip
gE5HEYFj5acG2krDGHbrL1KrQP1oBCXi09vWHVVEmhWV1WcmxtO6Ni9DTuBNLqRL7/K/DeQwtneu
ou8Q3clQLNAPmpVQRAVQKTOEAuIWEB2emCepcUDLA32i3ziBXUhHGKPpBVz/yWgGeNMUdggYH35F
toljMN93ASnjiFDh76K+MDixqyFUz2fCEwTm2iWmUU1hU04sj7mh4TUa3q0sWsQcT7rgquy0ei41
GO4/kDVFc9Qy7U7G2eyNPYW8q0CwfsqbYFjgu6NtVulMDHsEBr/wNWLZ/0Mi7TrVP3JAyynw/KQf
4N4PezWkjFSATS/Vy97sYoy8DHCZNeXmtRqSkif5IVwACZxusCBPg41oEzQ4vg/R3Iiy4Yy2zLQg
qChQPngYpS+STIUVBtV3zQKUeMCLeKfx9MP2ucyT30mICyQvCFyESw/EOqJDLSPw8CzxP5XKVsrp
V/Nzsbn3VtMaApxYNfVfjV5YW2mDWsA61PQbwGL9Eq0Mcr8VGnjpRkplUOJ/IojHsq7FfbodjOn2
0F5nuSghogrSjpgJEftwhSAALuRVBi12Ea9fqABpE5fIY8570R5f1n9Tqy0tNUjtbmZNH8PC47MD
eSDe6OUMNuv3yuPlF2UUOyjJuuiJnYAe4luLDwHjaJmkycYISZ2skCLCxHzuCGiI0q7Kz6Iuh/4n
AOjAvfU+r1rJeaxd9HLn7fS2p5lFcAxC+NEEH4Ezu9fPL9pzSz/KWx7tWi/YKlJpnC2fjeZiOYy0
mgT8sFDZ6ruRRFuZO5tXlKg+nbXwB+dYpH2n3DtkbYsHCbf1IV9nzuIK+D01VOUeaJEb5OPg6U6H
pk/Ala40jcUPB5wTC9CAqHKIHg0A/CaMSFI3QL1gnp4zXkd8prsuj5o69cNrPTwhJbMC6sjURSWm
fVMJlrqO/VwV4IHRHHKUAhznSlkqqN9Bl7Za5ek+YalywE6ECqvt96VHSjex7fkBdJOuikQL1UJ6
UVlCEfnmnMSH9k15FPR3F/GmfGNt9Pb8Il2HWFSMNvSmVvkRiHQnwPNhPh7krQwyX/cHAMq3aoP2
DZMtXZTy4Us81zPes0LamCLAHR9SDLCDAwCXwi2OhsoX8OsSgcXmKUFPTPa29NRaNQ2LY0mNoiaJ
tC6gTfwpgDGUe6Z0fzXaTYbECOtOiqRSeDOKrvbSh8VSTSvJPxUYGIvFjncTqWT8vVtmtBQR4cgz
2kngnoObl3fLiQpYFod/AleHpy4j5HRQALhT3e4EpSaXUsRrMPrE20uCgdxXLvqvUxhAufgj+7n7
KGZxzjDC1yWI/mXF62BLK3Cv2pPXbKlUa6ddo34DeImLf+zgsyA7Q7ViS3wHJ4Yaut0l/mq7bXpF
3n6wlL9PoNvZWNQgkaLeq4lHM1L+OtoSnOhTLkyOisGlqgwA3hG+sRZLffiY5X5KPI9mDA4hT9ch
lQIEvHwVZUYaPMIb8da52R19MUF8SVhxJzua5nQVLKFi+QAbt9goJSq5iPg3Pu6CIBEbz8TWTWh5
EwNRkH7q4tTZ/9ArVGmRgQ7mC2DDDwGs2cg5FA473U/r5mI/KM4mAYQMC/AbOvposrXYZ7uGsGHU
sgNrrHEvEIOjZm9a5guZopgog0o5CwOfp8Jh3AncrrMKEw/hhTbK2elwfo9bB+pEk4H98esHmAfQ
+kWnXczaRYr0IAbimZDUsI1JMoZgsd6c7GHcWQUMlMedgwb7o6u5Iwzsj7fq3owrc056eMCF26fF
pnOz+kWT25ZOAa2TjZOVrmdypDfHW8tn5TvGCtq3w93de5UYqre/RkhgqqJvOBheTvdJS6TqubNP
NHdw4kxmgh6+9mDBofb9pbvtIfMIcl6JMTafvGblo5CCWiQNvep3zh1teaD2E8RCJmhOj7n8zmwd
I74o63W2OIaWE+ialB9DSAI5s9HxcwvO01DMRIN3gp3T1f6LBz9/iAC4J+TEH6Rmo7uXqytX0dxk
AShj4ONQuOiQeC5Xr+IyMHIvnwtqvrsoR36aDkl9ZUKi5BBj9ytWi/4j0eNrzxUHbXbWNO7+Ev1Z
lvgzugPBhB7loZPjXEK4xfjpPKWlR3FBm23f25CmuP7V/hxpc+gqVBPlQTG1PDfUF9JmYoC4moJV
AQvTfrvf0ewGsab0shZfZxpfO6bwprC0lg4ZaoMWzZSfcMcV0eXJbYjgiEURoi7asSZWH6uZ7gC6
ZqZrlZm+oD4MK5ngJxcCXyFxUoPeJ6ZmS5n51BSzCzLXkYibnt55gAlwU1vuqTmV7BLeT561FMy4
F8tCz/QkrNfXqRjJgs+sw5nDSi3w/A8g6CXPjLkVN2l6huwNSxPgSwdO0Ma3raPvjVOgNsS5Pf63
u6187RLrBBaGTWBbuJY4dOUdgHLBVX++R2f3MvZBDtcVmtGgfo6G73ZevNXRHr5DiX/xoqjGgXYi
UFaeNLEFmtzhlPtM7qXGlaz0+A73GosPLvEthDZ5y0I47ucuQCBiQ0xHeKsj6CDjVN53n2MrH0xv
e85MeRLocgL7CcSgfBC35wqi8ZsjMnSA9E284ail/FynJA4rfssM/RXtte+K329LBkFqL4H+ghTt
4/ynKVO0lQIKIlC/CarH6xslyRPpk0Kv6IKzOEb520wb0SvArZn7Y4zTI80jt+01amL0fUEMMY5D
Xm4ZD1Sd90g3Am4Z+LMoiaeATAdZPDvSk04+EMNWEmLrXuz8qNjbgzqNFxUwqpXJZvnD6FqDZ2Aw
8wYK1GtWGhDwlAlT1oOQDZINa1ndR10iOh2+KpL0is6+8YhUMmfzTASBLHLqx1RZhxgehpHaFgfi
nUgTz4yNEvUPqIIJ0PEe5BYkKE1qOTmRbqkj3uxrmc8AE+Dp6DINDutvwqYrE3gyQejCLoxE4txE
qpPVrSz8l3l0xMaxQubbpPs8vjSXJIHlXj8o552y1AkogyhsFPF2g+dDgvT7D8hODcnFip+1bgSA
zayfTZyEtsYG7NvJvUm+q8hlPTWGt3ioRZobY3xZe+Gcp5vGF5D49qgzzWxq4bZduvyu7UAxfV3f
ygNgLUxlHK/LFNbf+u7LSluQ0SCZ5tzsh8ZGbtG26nf6+8fRt3HdnO+gi4zepnb9KDRhiSsLMLki
StPwlZIYK7AmoheJL7eBZeWdoNnFWL/cXIdYc6Ho5gWMy0IFfwil04c4wbunC1FEK6i0qugpaGAS
CEH6MS2qr6c7FNJ5Px7iYkH25JoPp/prMXdVXrMA0+BDryiEQoCpdo6sTLWFZbCJyLNaA0fBwzni
89V/unuLoMkeRaU1+m3KyTqMjyCIXDpm5Q+Vd0iifUH3Ezc3xDbVStBq8hb5gP1UPh1MpDGOe6Lu
wMyFsBDZ0FjRmvuC7hSg6M+hiGHtsEqW+u1bmIunrfmxwK14C+CsNEz4H+LBJvleuuKQIRz+HYJi
KXKgBRdNWEaAT75L05YiAwtRMiAsaZHFNl6EBNbeDdxgdCXrrM0TpX5HZ3ergDdWB4h5QPE1PcJ6
R5SiCTbo6PQC5Z1YpkI4RWPgX8GQU14E5mcDolPfvU9ZOuBlc7YADAbU08hBNYN4e6Vgg2+2jSzx
ZtskHsmuP1E5m7zTDaoUom9gNnbDRvwqhm/aMOxxQi9vdOpYzZNBv4TInCNjSz9wH5jZ/oyx6gIJ
qXUtmJ/gdneD+klKMbCEuKQk2xHb4VY21t8NCaFQt7YfsSqpzdYFtaJmAP9cg7HIABKo8hUv8tco
oT+iEV3ho75DzfLSTrkDH2/LcAis1fUxWhF5dx12kUIFVQz4oLlvJUgqFgOu/Z+hhw31VnuzdCfO
2xh9HlbwwAt7AZOU4qJqqSELtZ0Vsz673nTHrPJslBFQXfhbs4A+lYiR1QjhnRkCDfCKeWI3wCXa
9xP8oPxbv1PCSz22eEeSH5VbUuzUwXropiwU3JMlKY8YkoEJ/YeHwG8fk3AYfiD1rxZF/gC21DEw
fik33DF89LefjQar6N68iqIGWDf3IxpjGUY02j/SXpXlLLyWPO9dkf8sWvIraSCX5JTqXUC1klx2
gcWn2u5uGOZLmAU/OXLVW61soOvapMCkbwtulkAynZZeOgXx2OidufYVvU1YiGBBFEirRvOykEYr
GjvV8HvYkSUbIT0K7du89ZzzE/9V7Vexvl2sErQbCBfdcrlcx4rwf0rrmbYykkqVR/eI1lNEsEdD
0taHmvEOz2DLcdf4fQMZBewJ6mX3eeZubfJuE8KHy0/2UC1JSL0BHhk/l3LRhexdCM8Jn5OIUV+Q
LDgyoMKS70VNbYMjTbOwVqzKcnPCKCg9WX8DpZLXFOyXEyEL3vjB8jhmudt1HE66Yx3BYlnn00ku
2NqWbhvAQLqs5R6cqNngwdT/fhSFILA+TBn5JuWcu7BZo8giprEFaKBoK2Wtv7528nfSfM4SND6O
U1EOt6AGVbAYLE8KcFiVGp3pwJzCx2ZXw/uhUaKkeaZNnO77rk9382mK+4EhIMFFTNo6GdALgVyP
2ICcDADUHTcfL4RgRHc7DdNcOZZN7s1nufdFpS0cWzxGUhkrPis3KH0FX75623ef2ocoJ06A+hG5
sZF1HMbBJdR8sBrY4yT5dAz/aqUUUjfTGH4XnmodbD2Z8AhPIEtCHrr3qWFmjMBauav2zeTZdr08
o2kxrum2sMaOT/a4EY3dunUKxDd1EIeuVjSyULw6QdW52b8WH/d4K0dELx668qPbJCEmIfAcXnhs
VYcm8Mv22VBiCWpB4ODW30L+8sOabvUKiRzt4U9lKRPBppohBxoMUU3DDVGQGVC0J92WB+Edo5eg
/D5s8thLLh5msBdlulKDpR10t9pSnhnx4BGFbQudHdqSVwnnR3Uo1wlMVCUrLDOQ0goKIL1QBm0S
cwM01W0xyErjzvbdfs8n7Uw3F//z6TtcTtXMHgZUDwk6qzJHOtAjdy4Zq2gTRA6dFo2HVt+Hp78F
KYK9rOasYUxJueolgj+zyI2NSBjOSGaIPi76RB16gsRGl3aa5gtbbIDlzKT2UntvtZPT/j2117IU
UPsYiWUjQOHO6MyyP0seLuq6qaa5pLAobEmuGBlYVucKnLnv6GMoyFGmTU2YrX1to2iNDMpT7SYK
2NP5y19bXS1Wbb6Q4EXbnlUHUDW3Vjh34o1x6gye1OExWrIwNz3FcASrgcq8XY42M3kI/JmBdsf/
zHyGSecqMl1ii2ia6K4DILUyUuiVo0RyAtS2hjxXSNhTwnudKqdB6/W/+hK734KhNzjzBg3ZMT70
QbUK6ZxcPXMANjrod+XgvmrP6S83HJaxzqGr5ijHyT/LFnIZuD+hvdynJDUGPDyKf7WBtyyLbI+F
Sq6WD+XyKoOt8ltPK8WaTneo/dwMCQqzVo0iDf8jmDYfI9C4Cc3gRfvgJRP42GEVKkzxFxrhqoAJ
WKy9aXJOy59fAuTKqeUwTqKU46jxwXTk9098pkEHnc3rITLUiyVZa6VbuBCPaw8nKFV4XYzAWdtX
OeuruxQqdzR3Q3vmU8HxXE1ZRsE2yFtlunVIDPxGiN8WD9eCsiOhamPGeJ+rK2nv0VsfqhP+Ep44
UULVegF9Dli06js+xBaGBtjyoGwBYT9mOOEo8klwYSWu2g+kfNjCYxruJUOREZ4/yR2Ou1q4F3/a
zD8UAVhFPV5JeQN13tdBmlvsAejv2SJVWh3LgiXTw6hEhwpSxdjEfuxDCYhqriX5Cy/BiySBolKr
dSp2EFIO/H/ch523iBv2LeBtrhycbPm/eP6lZom+PqQsjhBPEZqoB+/m7jtOVcVv+ri4alc1GESa
jDBoUZcCbkz8c8+wCLTaBlhy4EzbdIpuAWnfLoaqg4vP4vU7tGN0sjA48MJqahrrolEzmZWlKDGz
TKqFK6OF1E6btsUA+yUnGYF4V1EFBq74jyPU4cUgYDmjFivH/y8+daQW2ytD9qOWPPJH0kk4z5xK
cJW1ax6UHSay6WhXTxjALdCqZEFBl3fXE47n2Du7PgAzpRFzDup48K2bdHBnag1g+oY/Asjx9iDF
t6iKo6oNpgiuG+gR/X4JPHe0g0EHejsF8Ej9PW5+14VUh2Yvc/CqXLboUi8wurnp2QWqFt2vaEc6
oKNCt2AGPIBE1OEcgZ3TbYvPggbyJsf7Ptv0deZpzYywGpAjiAIxEL64Wz2brT6Vhq0bpEVY2ogF
kL6+EuNdTO8b5Dx1yF6TNEPWYr9NWtfRKDucYrNjwqwk9wTuOrwiyvIBefrM+d88bmECLWTJ8a8G
s8N9m7MFrAnIzHI8AqO7OqdQ70wK+lj1iLqXNHBQFM4KojG84ggCSxwWAkcxDTYA4ftdSVqmAImh
AOeUvSPCBu7Nyfg8nze9FANdREK9y0MHJjElEARSHwuttVnJ3uV73qAG0NUSDFPg6zZwz1RT/KyR
aBXtHMVZMTJoI3jV90QBoFt9ca0c07QxAKPMnxRYsNHvpVtsgIEVSv8En+ybubOERbiRtlJOZ33g
pKSuy77FxKmsdqYFLLGQrKqsi35kEfRCGZBQDOquWos0mFsed72I90H2LABrsM4/ROAO49dfe5iX
MP1QEzwUxRhLPZUPAIM6nIpJqlNh4n4K137N9kmC/Tuu14a4kL6vlf5Zz1WfE6MfNxJgc5NgF4iL
1zQ7/loG0RWH3+MlBuCo86fXIE/dEnRL1CyMjmGqW9Y8xnb0f61Z3KbtqV8EnOfQT6xMJGg3ACoD
EOUluCOj/vFB73yOaoFLY/gMh+1Z+JvOvdHUdJcBd+7TBJFe4+8rug8YxcWl18S5y64Go/HG/s51
rMxFT3q+oVZZ1bTiG2TOpzHSyeL9ecdl/D8ZoB8xIUFOj6K1eVIrmR7SBXJtuXKYDJKfdo8RHC0i
cxSVpmmUCN9wK0YGFtf1Rps7Eis4p9wAt7BXIRw/A5OgddhsBzbIuK+bDpfxCoDqD+rQepKAJWLE
j3UCs8yr8K2qzSEFWeM5XOLc92wkc6zS1CvdKOzPnrEDbCTWsfpn0qUpKvIMoj+VAkBgDGOw/04Y
mU7sT0l7Z0FOuPEzCW7PlqCX3tglYMBcd3B2T4x8AbUWvOSHiRmGTIlhV5NQW7LkdmL3Ej7X5muh
X3gCKviup5m8zFR70TPtlQgew9OuAY83cgF47SZubiHL1FgkTm6VRbfQK+ZlhlpA6WRxJrsZP6TD
WBDl+MGh8jQODNijPU9hMLcZkDPR7yErhQnUx3U/tiEsPCELpMT7i449TCeLRl/KwxM6s773yPPF
o+ZutdjKRqY192w4m0chsk57+eYtFOGMQb5vP2WT2Z3ImwYTWMBHfOf8XwpFAAbgIqBfobKY+ZsB
f/rQhfZp9QH9J4cJkr6VkDTNFuWwnAYXIsmUaP92bx/wAnu5plT//m/AAe9ZDeXRA7ql4aIexEk7
hvymElGJlXtIL8F4P1i0dx4hpJLa0GVgV6bQFZsmHoHI0NAgv5o9DNjpACfQbADSWxNPhPj0bu3T
RpyFYSXcxn+4Cy/GPEU2yKXYz1ZRCm6ryv3r2oyopedTF6OoVOMb81ovHnCuPWmN8zFBpWpe9B2C
WDBttDiZqQlq/FXZ2TDoU380pkjzdaex1QS3DbkxS9a3L9msYDPDzwaG7gML+zW/sqi/rLQWrAGW
awhEXfezuPRmvrXiD7r6D6wsJJvLUDxD1I2/Oy0a6H1QLnFpSAwjlIxbuhhxiFKEC4Tol8MI5CIp
qzKG25yLdV8rGmdn0d8Mjuqzpx/Htx7q5AcCQksslemjvgMEWcT5NBSLdlk9Dxw0oC8oQAD3D0QX
DCT6K6W/FImeJdui/7kK2VIgCGxMRtu1w4g7j/7fInMCo+hbUrJ6VoAoRd+6aUmLL/X3L+LAa2/n
t63Q0++dG+puEU8hAu4t+NuDsL7veRkiRV9zhbcs6WNQYqvl0C4oecfikBNkX093ijmKk8aM/Yvc
flE9jTHuCfUGrv/XZ2ETbOjl2cwfSsbmx9qt52wmgf56xtfEEBcoqmYLfCaCYltJXZ8jfV0X/Q52
K9j6C+GRSJ0HDtaavtomY2ZOwUWZ6HZrdNP8YwmJIwJH4NXnY3lN6ZF12oD64BwGw0PNacjYGqrT
PAgiq3gq7j2ohaHQtl500kqixXm95XN0qElS9xdde9KoE7D6SfSWGyw+vmBN50zKPmC7domP7btz
Z0hu1yU2tb8otQG7LZLysBZ/8OuAM9QaH4WFyoPjuNHALDbepvuWC7JWoNpSudW+sxzjYiumYhXL
u6CROaxw9Zq6SqrZ9nMEyvesv7SMJoRigmK2RjOuivNgwUcmICEfcrvi8J8kS1WIVJSF7yvQYBIR
27zICJehbE7PoeKms1qZmt3FkZqexR1XeCUjKdOOiaviKcgsEnE8/NyIBBTbty7/tjr8DQxHQFLd
ju4PF9n1gqQEmVUKui653rA7MbdPaQQgqTP0XtvNQceNyFXSy1b4nCPqvxMmFeBrGuCw+FsR5Qrs
42KojeDTSMJztymP+nhAfvLAIwOJ/0DQ+MjjNamXkhC+PLmjb8q/fvP9JQ9mxndTSBqYHg/zLG67
fhWOwRWyaPkgY5OxgDEYp7iuhw4x2Z9Dv47rwGZSdPk8pumxDGFpH15nV94tOJFiEEplfHz2w/QE
lS4UTOforuNCVi7lV5K8UJTqxMFRn4zW3CLnHyfjizMCbUb62nVcWqsfmVxRBY/RXjiTKJmEhuBw
EX3l1PW02RRKEhL077Jvi/p9Wmd9ZflHZ372smYTv7nwqoY4nMlWdDOnyqpkIiMqZGRu3ovfaPfU
de8xW79xGUGF8rScOGMRkFz2q6ZkA/veIt8Esbd+lcuOcN+WkndfX3V0daNhVuMzUJRSgEq6KcKK
B1/hmQI8NKxQUWGFVY3Ce9dmravLYtYu8R69qiXQwADCJueo7QzEDjFm5I5Rs2b7wC9K1roZ3Qzx
w2xWz9K0XM0/tIUKUpyOckmgIqmbKuudbY/v0F4+ANQ7rd2KMnM9Xn/epRPucILSGmxUvaIIGWWf
ScThVkh07p7uAn6rB7SAi+5VhG1db1vE3U5OdlP4J2oFe50UkBP7x2vYKLenu7yKDZ6CuDJnqWiG
VTLiap2uhymIElXH61+kQCIS3wI9jnX9IzXXOOqn06dG+WVGgaGaL20hGyY9Kmt/G5whO4N5tDL4
ROSvomJUCtsWh3sXrnwNBsfF1zUD2oWy7xEGg2fPEH4uFjUWdTGkcG4xCz4bdPyb1P5p/nfYz91D
Uu5Xqwsj1N9TS83LYwn1c/BJyLcEUCGpdER8H1ZpDaDEtvgj3sKtKw9ZXULd5178MAQEtDNbGvwk
+2GGr8o83QTQXSRX/hXv5o8lug/D6nsQAunr1NN/gINmTur+Qr3BBrUGUkAYysBLaTubGeI9bBkq
lTbACrimkyo+wdN/vS3S+ppGMPt7bgIistLYx1XHxreI6HkwzQjH9V9/HP8XkFlouo2/OHHeN9Q1
47xY+ioG0qdOKXIv569nAnTyw1A5MWVdGzwPjawrXrAcMLpiQ3LmZQvlXeLT5+GgZqrnLzljcAFk
x2xc0RN+bOYAZIlVmItTsH+WGQPspFADW7Qp36qLRi5Nu9EYa2VuLjVARI5GntdEHQAeiyp7Flrj
r7SPrdFJwf1OWb/kGIhZca9jwsgwb2QXUwQdhHdL92Iw6FRnDsITZImSqVl6s/w3SJRi7Hhjvp5c
UdwFO/eWSbDB3WsgqPp/or7GwR0ZMb/EYBhTNzOhCknrhyvYXRAalTkqixHkXqM4SsFUNWaD8h7V
++NNwhWAuKtRW1ymOjPbG+hJO9zCsakgHTEfygmYDZhtcPxLzhY2zsWiN7OW3Xdde/Bm3a8y2lid
qFHbDKTrUV251/D0g0OiUkYEz6A9NCksYe3FqqTcje/WkQWhTipg4d8TKD0hSQMPXD45yg8zPGoo
xB6e4OvDmykXKmIHZ9Yw1dNu/D+Gx9R2uteAqLsvNiztZuHZRK1xbwEidn0DNAhphyyqVFbpgtUu
CwOGZOyAjCJQhTd/6y+qF91apZuBr/3TexJIPNu3eD+8ua/v04rEzcAEoAQW2eB0ikfsIF3XVuQA
789GrKORqUhEfT4Enjs53AwLU0w3lB3IED8XmCeZ63rQIRmmrZEcDc/vQQybhcI9c8dKrNuU5Tzz
Ga1+dUZBDYMRogZujLn5AamYYmL/ILia80qecOXErRhc8uRAKX2s93Gf/CfZKT0JET1SHibXdbo8
lsb4QTHmvNwUlPAeUza7F8KMxOe0Y3W8noUDBamyMjMd+b4TCCnilnKpiTiOt1EqIV9anwLILGtd
R1povNWSYth3V2cRHQ0OKb0GUAQF+jjArot2FTFDaeyM+1kFpjIk0AAJzI5A2w76CQ/e+4JtquyB
S6L2eE964SAEtgFgKMAG7NcgrKUgQhQGn5fXTiSBKlHI7XomiQW8YeL9N0+5FKnGxiLirA772Cl3
1D2NXlfMJXjNpEoeUdLShc6hqZaEVMVP6bYHYF7FV0xGYliwpzaRypsljVS6HQYtNZ818DRzlgq1
LObMP66c6W9rg4eqnC/x8TVcTmesrYO+aryjE3gVHohZQEhj8/ZH4WGNrE4AKOv3rcwRk15SDEbs
rJxNFL7YpF+wqExHHwIhk/xKhV0RKYO0AoRP0f2s+dRQ4EtZZzE/sDhx7UrYmtcap9zObCQMYOee
pK1eFkCA0cPpgD7/hXtHeXxSEqK9Mv6BRa28xOPCr1BNNdyiN3F8wPIkkmSm1WSzwJ8WjSmtVOg3
4oonSBEAfULeoCv3JT3uIBbLLNCdbhWX3wlpznr19/UMLZJL/UluzBRAQLTa9iJhsHXNnYuBrUYo
RoAtoWXAn5KcuFgtSKkoiYa3TPVMiJtbdjR70V9dulXqp88SKkyZ61BviisRRLskZz3YqhHc0/fq
XoNKjfR+XNIZH7fH0RDZ88snt49w3JPH29EfTy8882wSbSOF6+JyzkMv3TKif6bnkvGs6OzdUWvd
0Yanf652rRrcVeHnmkGeoUT6LNf60n8FAe+Tk9vqMutSip+X6wg98cR1AuyrL45Ak3PJmcd3yHrs
pif65CmBHQcoi8KMyBYP6IPzN1NuMv7X4vmuXcNv0d5/w5Fz1BAfyZwnJlpCjZbc1YHYATQw9HGs
NWvSEyu0pPiwX6QDLzaoXrzK/5hX+IC0Il8iZ/sCSbeidL8n9ZdxNmFryOP4yQRcFZ6N4oZ4TT7e
EG/96Khie9YYfKO5ZLiKkIno0NUYRUIPHxoFrfUrtPl+vWrl4lwgp61F357UY2uOOQcNTUmPwQY2
0FixQcnu7LlMifmOJfL3wFijxccf1oEDHn4WHwEpc+61LzbrFmMryiPddjxf+nPP8q7FOGXLdaka
hs0XJWz85Osx0JDdm1XgWjISea/YApOFEuDW3m0hveQMAYVDoKGM0EKnW5BB2FiPtdazrOsqd7PJ
d3AGI733ciB6Cj6n2uRk3n2YmEga2lKHTerBVA/b4W0qQAuZMrFF8BFdE+HTBbp7DZVtOMtKReju
XaHX0TPSA/iSMYZWEcHdXYsEuAWqFM+zPLcekESL5DmswQZE6bPMLpzIHd/Sd90zBr0ahSVRtvv1
xQQ6EXGPdAJgBFmNFhcqu+h6ecJiOMEwmZxIs+6V+qlT6tLpYomCFVrx/xhbl9YEHWHBaUnhwr6I
Et+VL4usbnefnfoHK8yz5Z/NyKVbVMwYGX9kaSBUgGCEAOEOF/7/IkMAqEsGVzZ1560n27uHnQOW
affD0yD6ThJUbt383WXThggSJ7ryqoyOuxxMv0kF9UyQzL3GAccWf/8GVHfKaOFcuomgxOKD9buY
NepbXMCJQxMpK+TlFHee3v633+Pztb45n30nJ01JG212cPs6/N/bVUjXP3iNP+e3+N0iux+dTdzU
C+Ddlpo2pjgxUvelWPn/rHTxzyeRbmPHt6J5JufaMTs/uuZWA1HuZuXCxrnHn1zneX8iZFA7mYce
sGp8eBig+B78jFcgS6/7SZzXq+9u3q3xkkT00s3SImJFOTL7fNitT7tguhiPojuzbAUScrtgi7Gh
Sghgt0kD5VN6YVktY9JeSqfCtyMGG2Z0n2orK1ZoM8Z1iX/r+7vt8M9YBLOmxS8R6Xmwg8BX39aB
iIHgTJfgHaMPfe1eNACaNnzOMViThDAd3vSiHiiPovFlu5V05hRX6hIZt/CvjlVcg5BsDNCsK1w3
DwlJUEZh+ADt+OXlzugXNHQoVqouuF7oCdoQEWuxZI61pSZB0fqVP/zOcY8Bh9FHpAR1lrFJvmVx
NUkuyCCuo7pwiZnUJzjbVnW5vom479efLBI8e3McF0FO2C2i+S5DOotHUh0E/aOAtldDAwcQvG54
b8AtCGpShE/qx6sVNXqLDJeaJqHqZakaKzuplzmqpUJ6dnSxr7sh66HZdeqewKWdaZabOZXCqzMl
yyKJtKL6QBq6QXDwMtusNTF/GC3Q58jWg1CApaZ/UErYFcm2v+eZKRpbQ3fxTGcmbGtgs9UJ4Fkx
ywS5MvnV27FKSMjElSpEENyPhnP8/ugAM2Ku/S4bswtvHGbY7fwZRkqiQAP2XICzzC1BqNAzD7ka
cXUXHrRM2RxGwFtQiXm8IQ08l179pc9yAGQeDijzmm4Nost6nMDZoudCKIf4TU5qgCAd/vijvDV3
O71SoJVACWdfSWH5USUrIqKen9DVd9NMAMqN3LeQxWqc/jPxLoMUu7z3OVLF/k5U82893gpfxx8T
Ql6u02WEfSeQ+TXvXqk61WInW4pLUyOeHpXJXMPGqwiD4EKN1J4jfYxaVT9Z/3K4q/znzs2xKZw+
/9tn3Y+idGcfe3x8136+H3lDvcurtRzT901ofHW3V4Pr/8Pwo2eJyScVstPAEjpKvWPi3Uex/rmB
FY0BZcpyLASWsJXMPsjyHGxU8tttgX46LXZv9y5SO0vNTfZBa1C8ty2gjstkJXLKz0Ty3/qkw8QV
ZbXypMQeE0++ULHYVrYKeyYfq5KzGklyHDY33bxvaeKePu+XI8DamD9UyzDpf2DcLLOhTk9xeoRK
QdLwwF5SOdziaJt1eNvLG55hWR3FbHzv3AAAtf+y9gcjuKWXJRiKOry0voT1yIvBqBFw5yrICJbt
frQVC1FPjM4BPFh+H6Iqugdlku1bY+eKwKw3V2V8W6wX24U8/J2b02OXglXDTdrB3ToJ2XxLTyj9
xK7yrEXK2sQunacm+VViPNtKJOy31WgTb5Dw7hq4fl48n6xm2pIF1YqXrARcjndBytu9peUqnfja
LwttwVmcTMPvhOUDItFMUuJxIz7ATYzHj+t7NU7Z3uk0qIxyAZjmlChVJnJeXORo1zUHpQjqMYsu
D5B6Zk7xOBYrDjB5yrJ+UYQ7tS6J/0T3ymRjB0uUAVpEkjTsvETzQYIepdNQpZmWYGlmyiuISvIt
WJqRxAKzcEj0QTwnW/AG+sPwTUoDpcOe4dAoc3JQaK4ORhP3zJM4sTc3MQ+214F7kdIvzQPiuzZ9
XjgfCyaGhEvil5m2x7m1m0u1zvQSVqiKBQNh4onFH68sB3YDHBTdHPC5OQ9e7ngfkopexI1azCxg
hm5yGUpVz8zzEGV6Owj2NinB87VeNnQmg6vhpwsOZB4XnCz8F0o2lHa3MUMWekGz+/+xJ3H0ULF7
mhvwS56oQp1/OSlUoNr8Cmb2wC35vAnef9Vjmc1mfAZF+LBPUZ8WVQmdqPzOHXlbeMNiSouyIbdJ
SQ12mPLJ/+X+LLlqA1q2oKtOW6chM5S1NP3RVXDfW9JAcd7sEMseviacOYFiOwKCH93gHI6xMIce
PWEca6Gk1+gXq6zeu24f7rWFIgNoI01V8bnlcq1/g2inYOSKiVt45PTavnup88Hbxfjv726QZGD2
0R1WkyMaC8Lq7g6ktQItSZQBpBN9pa+1b/HJlNuKsn8i3VmcxNsDyswmegJZVywgip/ere8/rg35
39+MM2nX7fJUxde99XEUGmsVzoXjfGknG8Lx4chm/fVhytZgMGFHjwZZXHndBWRrRTqg7/8N1h6f
BnLv/hiuyM2VmXC2k9WjyhE+anjFQHp1VcYYpA1y5+7cCPXjxKNlIiHFubPuzfl0B+cra/WV1Q6x
+ld5Np7dnL8T7wZCir1tGq3HGYVfroKLtNKhbRR/FuzVzvXW+ZbE6mjj2TUjc9DMQUsCCFf2qPUy
XiVcHTzU6H0aY5v0OitfXcRmJqTbzd6gTHGIYYSBDDHnjVY1w+3YA5IsANJQQpm4ZKu/F5GwyxYi
s+xUqXvBFaCfVY0mQSzYVEJw9ZvJ2HU6Oicc7t81FPYMFcdSxYkqB0+hu4kYkcJSmiWxiVh+0FO4
s+7iFTuEqlX8VPOliO2zabPeaG4SBsc+qQDEonuJEdHQ7HDfuEzngoPK7NWBkiiu4b1V98eQsu7w
MVAM1GWfpAYrI/so95jGuBz/355QQBMljfNOclalpeVkc16F3rIclADZl9n7eZoAO7dlWqw8gl3H
7LW+w0Au5N1ov7MK9zoWNT/g1Hz/8/KRwOnq2uiIVTyDeap4CPFG89HNV/wg0PYX9lPuXHgX7JOB
dwPCGJUo+BpVpvWBEEq7H69hJFRDlhRrgaSc6ah9vDKdjQW9EAxcFi2oA33aVESGZu+7vSIp6sBo
Re2MPeufMDqlIRiSw+gZ2lWSrXmWBg0eNTnYXg7dEc2mRGJkT18yHJthHI3k5KBTZYYooC/EJGfD
uMdggImJ1nHrM7Dfspzs5Vy/TFpPpNO4hsyRslGsxUS34Sgavg/v4XXdemob8LrC3QUN49vDB0O+
mSf5B3X44SkQgp5TAZsUI5dxmdr5rWo7/gnAbYQeyyTKlmjbEtFdiTYnGjxkTHG8XuoGMIQ5IFQQ
hF5E/yIQMFTphYq6mW+wiNaRxzeRsF3IVmaNhE8QL8mLOlsaLDzeHwXSmbN+tXFuEz1bC3dRLj6H
Pgx2FbiK0fagEbGBAxWF5Fbaw2W+1yMZ+NHR8fiDkHLQbn2KicnmZs9wMs9wqGL08loUlBhuxfn0
L4lQYGMzUtuMPbHQ643KJxc2B6W07cYRxloMEgmcRYkWcS411MLypSgx25D70ESI8Ya73ZptrAka
7CnIOdRswKYkIpD4bp/A5fSBlSwMzhLKk1iQEZiRxJVAfPfmLNPDID06OU4/+AsWyq4rMjgTxq1C
LlW78UVZZWqQ8tikAjV6/bvoQK5tFMV0I8VXSmSLJw9NAUQpVQiZoLfYxxLnH4XJKvuYZ3YibWmv
bAj1lwQ0if0ISOqyQqoPzfUNvzhEtx9cXXhmFUI4R3hZ+IkK8yrHrkE2qRArCUKPK9tobXKEqs0f
3Ef9RE827HBukKd2bJMvKWyxZuO9ai+h5Qf6eclbq55Q6sJnlfpWq09IOK7nIN1bfugn7slx1QMg
g2Gp/hHQdZ0ZpiyBGDZqZQjGoPnNkw02ChZhk6fHcwr/oNgqwFVaqLT3K25WjEB+Pr/WkVeBL0Wg
Vo2gW2+nNUMlRgk6Sov9llroCaq7I7YIJlvLFkqULoegohxIT1m+P51DcUXbu73POkSm2+eNOSgC
+q/2jpCjvAeUDCMbA8SxFRwPGK29iRWJ7/lxnWpdlJWsVTeIfWWOM1mcB1Mm5+Hl0qxqJG27X5xt
pOfURJuat/SP6YbOWJvMhtQz3YVR6lNQbPu31Dx3fGcHgH23Yg1Ns5OKt7wKLwFQLM1qMmd8ONVm
cf2odccGLZfaePKGkFRRask+GADfBoB46/aEJWngsyjamgH6GVQLUKs06IBvetqewzo7V82CD3Ka
Tq19+WW33H7obGCqAitsWZ6t0ytB99cTI326I8QRrAFkYMKg+p2miWU5NhNQTJ9beLdFFM6zwtha
C1RPXcB7bsj1IisaddknmImWwB9WLvQycWdZ5mPkb02/m/k7/W4Lpm71ivFUZVT2Bbu+RvcDcBw7
DLuql4SfYX54LVKFN6nAwJlTKNmK5iAgKEb96hKxn9yL7/ZvXsQ8gFEh4Yj6Ebj/hwAsk2Hdw6C5
hIKP08gBXEtXhMa9WGXE1YOr0RW6EaJ0lpm42PavEasscfJOettofWnqhLFCOj25VmSpF7qd3kNN
Hn9/NkIoHCiSEn+7YegBlKo+F4NYtvoHkBrBVb1ZcQh1Og7itqM2Y6bYZbwuP84BfkQDnVLFfL/V
WCfZ8D+sb88yeWoskTsLhKG4u37wP+C1P2B13xSe1kyHSUQMsd4z5+e88EdIZiVHZSS6DcIeOqNB
PDvTMCukVlZpOijYCb0GNHGaxTYg7rZ0PKAlPpPzCmp50KHNCe9IfrXsSEjcQA83X/idaeY9+t1w
7ktyx+HYktJnbHLrdLWl4FeMKoFOLWntuCKSeV4y2rNyOQRC83M+80xSCOt/uIS9cuKkJa1LAyhn
LGdGMQN7MzCu3mXJKdy3UDQ+7coSly5UCZv8PywTyQlK0dVsDmpONT6ZvtGRO4Jblwj6AHlBpgbg
2Xknh/V3tc79VzXsGGfTmb4Kb4/NffGHLtOkZ22GqAKDh+xkT1OkSgZqu4KdnSOJ+HB8UGVgsU3T
mP5/9PrLAmgPMCbLZCkT81VEUf12cYbZdT5vZ3j+7Dpb9HYtB92NiLC6tMLnVfYeEQv8tmvtW7uc
LV38GtwzzxeX7rIhJWxX8ipTf3CstqHgudKHOT9PruQRhuNtVTCTQSW7Xpx0rpjG82sbsEfeM29d
cjVSpk7363JANtULAKyc6o/MlYAbihmd3vETk34i8tCWA5ijgOSJi9nKs36K5XuxJbGkVtLpS8ia
nuVpdmCjbG1XssDNtiq71RRarAiOmTV81bhxu0aSwEkq5I0w7MFuRCG6JpruyL4dncU8aYjBXxkK
/mTkmdLSrvlUozRGgmrjFPGxFfDrfAarYK73zfDG/71OgLSi0t0tIfXofujCglbM0W8ySGymjPXR
gcyl4x38vABT+qIgPpyUWiD2WiDHEijsB9+JpWeJwEGgsRJ8O05+mUoIKwPoQT9hSvRbAiKinW0Q
ALd+g6KgdBk0e687jmmVl80q4hRlDNezmKLBs0Z8SKpjr1aZOhLQRJUedgy0VO5vXZ3kMyPZLfJa
IkNV0lEZ0Lq70UXujFOr+hLYR6IJ5KWia5CXszmt/DufzeHcD0A/nwnZ3vV9RQdVStmu9KD79b4T
r4mm4e2oMIBVpp66JQ9jmDblcdi/d/5Gd3b4zmYlMg0zgg0T2jmIKjOOW5byFXU8U/rzeArBEZ1N
1U5fBm4qyTbgM7fZPvXP+Wfx7ydKkl6/3dPookD3rCwpJK7Sl/koSK0815hm/rZcWNBHsB7zWPp5
XIbYBTh2YPcpTASDgvkY+aWuIPRjzkdW92onqW0gi6lxw6M3JRy5I6v7K2l1D7rW7hnWJmpi+on4
Nrmt9IBs9ctLiMUmIDmomhjtrP0GUMDZ3gTe3GZ4LhD3oRmgYkZTejFo2Evwe2ZN4MqeGFPJRgRx
PG73R8l1TBJCasEd1ITaC+AnXsxBjD1S7DPcGspreu3HfrygaPI2s58gBmcWeoz5kCrzR504CkzX
kfnYh/GywLoETIDOf+6LyXfqUqvHDxzEx6VL5zuRi2WoEQcyfOqzSf7arHNeTeSqnIsDv5wZsHUg
D12x1WsNwB2cvFwj5d2nEDB78qcCRNjjpb4iT+R2LXes3/RQ8Hu7x9PhCeEpc3hp++pI5NOS381h
kJOB45atF694oeWULcBHmYtl3hxrrgJdE4QpTzgJU6JiWid70HZghCGXrxqkpyd0+WPtVx3VYPUq
v7dAgEaG9MyFUATNcb4NRCaKQKqdUQ/TddZ8lHVVldCwJebWUKhG2P0wGylrmO45Z3LI2FNaEjyn
POyg+fKFd6bALYsCOxOsfgmkGPHPEOOt35HKeScddsNmY7B6KvTw4QAk8Nj3N1lhcAcXFdW3HYwp
d2G5CiQyKDA8jdto2FfmRBwuRw8aPj4Et2sdQZs7lE3Trgy2Y+937+BljoMvcdoLOBs6TH02D9ls
rTTdnjMNfQW2TPt4x4o2IyKCE89qeqg3CFFigLzgIzcFSkg99orr3zlCRUzAJXXS2qrz7FgjiRqZ
EgSOlnJcFP5zmaPp3hHHW7nkCMohHzbUXBfNmu3A0xzKRvfBkNXHD5BndPZ4MXBkSLC6rVtY8lm+
0O4piEcnytm1/HLICXDetGBv02IEAj7BfSwYh22tvkWA29oZ4VnTjH4u3+nncEzP78+oBbFo/T52
CMHUpXV6KACs91HrNOI65fs5HZJReudcauFdedp5dWBOuKzK7KGBCz/ZMpls/4V7E47/ATNvqziD
ydKxxBWVenFgPM0uCyf+MMhqKvbh4CILo4fUwRlUS45NKW0icVtA8UwuYWqFQ1yvNcBvJy9vC7OK
8k90qlNeLnzsqlWWiC1McnZZ0OVUdK2i3tBUSeEPN5CfoWbfC9NMOk2PriYRfSvflCfY7+bwtdwI
f6JLbTUuu8JSqiahynSGF/9voMrlN8L9o22Xs7iXKVEgQAxALSMCwCb5SZVkXoMxqOxG1JANDZ9t
sLTrwT58aXL12BthwkXEPW93Zm14M4WYf+aeuN+Ii994KtnwAxsDDeWia2iHViPOoU6g+4RJ/jul
eugz9DscEw03PKSgA+8OpaZMNy0gVfWIG5OFVfa0Vlvc/rUBZevhzLLBc8/wwNmFFliUx1BrY00L
Z9SncEKD/U2k0Zb9+lL5IXTn6MN3r5fNF7CGOsDWFTyGfZGQsUkJbXQCofjjckM5SaBX+Xn+gREy
LTQzEqNqFNxnRwNngLmfGYHnp4JkoCld4IkW9Fkvh1flNzZ1ryKVvfSAz1VJMVM2u8ZtVfsLkhHI
BKE8yc3MU9ih9UlP//KUu4t46jje2/jn07t31ZF1FaDN7DVz4ziBbIJGtRAfy9sJCqa7gAvkuXFA
VCPt3Kld4/u8JiSQmeyE+c0r0dLCZOu0veumpShXv8L0KH+UEXMQ3/CtRSlgQWA8/3JgqGzLcbsu
3gfC96xBPf7jjo+I2wyxkqvC5wrR0KcLwaZPUd7XzM3EyXqR6FYYGOKHc/0wpkdAYx9qAl47knXM
OqKDihds40ZYTqzPinwZ0WSJJ1oMDdJ5jFpzvXropGc4dULFaEUx7S3eI4bXYpFlj53yOlFjG/mV
aiJnTgOj63IebMn7cQ/nstmdn7vNgJln8M5LzBcAOVWvvQsLMHk5LpeHwQ2f8b9Bd6w8mVCvmLvu
JlFikspkxXiTpuy30M2eKIyxLvvSHfs6wEvT6Joh91/BMhi9+6b8nXUTQBVI1ZskMrziVt14GRZ+
zlRO97SJsp6uCW3SroODz02Up3jmor0BChwZgJXnP4CusVJW2DQnNj93hauhUoMuZcfIpMF0f/Wk
WqtXGW48Ih41k7gK64ErUGTvslwhitQLpaZ23A0Ptog2nojsd6ZJV2wDMLctA2zb1RjUqHd261dm
YoO42xYw2FbwE1sEr7zPVtxRLcOlGSY86lAJdcrR4QDhbCYs9+2T5HOM13P5j9lhZn5NUY2fJaxe
leHJrOoVfqyRHfYCR5KgZbD1RCRZaVrLw353f5RX6a2qV2mndP4LLa+j4MqfeJ2vfuPHfbRXuYFu
+TvCDCGAZqx9vrOxbrHySvzycy5QhEDZwog4f1nG2l8my2h+uHxteod0+/JTqOsYS9ovLCX0OH1G
D7LAM5CUtLqyvcIY7XX0ZlzyNNqbs2lifg6bCMw08O84DhFDfixgoZDRa5LnnLXPkcIq9EA3OuLj
GDmCbSKCZ7Q8sYu5Qsac4X6WT4htVQK4VUSYd8ZydCXZz6iWFgmmM8FpAsv4fK0k4sRPuPQop2UN
e7glU2MFMymw8yTge2hhK6LnPLkLsQuqehiedwBak+b+hoHy4qmAzvqx/nQqdmXkyRJYhfKH+qLa
eOKviZ7Nq2TeRhHpIx+5QnKHPx1oWAP7S+iOLLEuHIjel58yESbIVwq5ThV+q/KCpOxyzlAa2h58
qUmtD9/lY11OPEZvFYJatxgIF9oqRxJDhLdA3skEukgZ+XHXJXxqBUcOA/VkeucRvSF642KyZ036
b9XrvDMnZcMUJWx5Bh2iC9m3ren9ljKoM1rz/eqN/OAuco+e0q4MI3GNYnEmOl38ylZwYs8deKVr
/Znp8bJlatNFZqFrFLEFREcBBw7fPY4eZKHos2iEDyg5QYZLB3fZyx7Qtco9UCZun+1Y9l50Wm9w
VLR8t1KUyeg7pm7Jte6OKNncWc+sU1u4shji2ArLKcWek2kLtjymdrJmmnGAr12epaFPWKCc5prR
m91H+j4e3RJyyBkwTMUzcvnx8rWUj2KxjnZ6PfH7L5Fe4QVJO47IsEPLooGWE5rII6Fes0dD98z2
fmNkJxHjsmy5bN++T2tQ6m4VgqqL3DcFcY6FfG9f9ISOtEdyudd0S7+BK7vYuyyH4+gNtj/Dpl2u
b43APWhi3GsVddYJreNK5b5bDIpK3HXOnyAjMA0k0xeFyeZF+sRdupaQb0zQn4HKzkl6kxgPM9R0
krDHsXLScT1U13DaE74+mcDD2CW0PGnnGw8QWiKeaaJDq4G30J+f0ERJFSVXFoHr5FcTEPmNK22B
2fUsttYh/2HL9bUv8YkBW9Ed+AEAoS0gngOpSpIxARPs0m7X93oCufh/MllWle4nDrNQAJJ6du4U
0ZuowALJ6nWJRwysoWBdtmydRD9v8rnvIUw8y54u7g+PJScPBO9+Onb30TfbWkVGmXXvl7wLEWne
wBIhCr2OA4ajrQx/p1CnCruwGC5FdiqmUMSYGxyjQ4xsvpD/e73mrUNkROAn4qyQ+T0wEhqD8KNT
BX+wxCSPDbz81AnHCbX7I63f5w3wUeSoxWxZbT3b6Aaqf7ytCwya+TnltBcbYHhv1+W+5MG6y/T8
Hs8ej7Q8t7r0bX3QFYqCbP8YKliNz+B2qYYP1kOs8GQt2DSaM2TYnXXsfXPZ3RIdDvQRji5z0G1B
VI4LYtJ2Wc83i+82ZGl7z7wBwhB+SpOF180EzH+aMXObuK3rV839HkegIoREUkD4DYelscoZiK6k
14bOyUE+2Ysxz0Dut/ku+PSzh/dzCMtPjsj5J7W9uNKIQFMw7Bb23odKKNb0a4U5ITcGumt6ebm9
0pjMtOgsZJh8f+Bi5/Dij1+fPNBCyDlfqe//NtD/bZKW7ZF0sPJq+bot33FMmlP6j2/kojGHZ9kF
74NPBiznXyFJ/+xcvZUA7bKuW/t7OkOjwOA5A5wUS69vx6xYfYX/UJzQqAhrYGUFXb1eK/lzYt89
DxUr7wcZ+ELUREht/4OLP8ytUkGXd4b3/B5wJ4OWl700AjIxXQxyj+j3Ptbs3LAYTD0C+w5f8sN/
hB3+XKeDPSFTCzwDnA6nHkcgX2df2D1t4whKqdIHnVm+PzO5izY4ab7vyEG/w184piEjsyVVrKcf
omHfLUoPTUQYrMGM1E3OgLdc/vRxtw19ompqVSggDWhACVibnFCTyjl5R4b7HMvrEZRUyxbE1njY
Yu6ROASzkpIquOTPkuxYFMudTzI+TK2272W2NRU1nEs8JCAUOJoUqqrIw9Hm4SVPmiKqnj5xqtaq
Stmdg161jcsFPamvvwZIQH8hxlHBihgn5KXNPiBkvBQGk1Axj5SKIOWgy4NzdvDHT/bk3TZLSuO5
sva0E02499MHR9tkU7ldwaoXxReaKj9vpuVOQLDSt9I9S+rVKP6zqNHdsAVGfpng+DmZfg0QiGkI
p2ODTEoWGnyxN3Pv5S0CB2OD+0fkq+EETANDqhGJ6Y1y0ZMCU/6j5XLSq/y7vaEM1PgoZVYt/LSV
mTBXVjj9ZStznxm3sla/bBBqJHQkxxCIRre9EGO6YKBD8W1FMsKeCH/mGLdb/EKR8KyVmBVZYV1R
IphX0Bd2C6Yvi8RUq4LeqCf82x+fzQcBw/goC1IIZC9/7H+3BeX8DRpbehnsbmjrAbP7+fgSNF68
3diY8g3f0GFYO796HubO+VbS7sZoJ/5jOgDiPg1gSOy047UX0KNcRxf3en5JVJkbFSig4LPV8pqt
ZG2Ba0bjNXJ2JbTMIaonTQngQb9Lun6xZ490KSkKllkrWtoGd4Gnlq7Hw9z9Z5QjCgsfBjaTz3Ry
vgtHGluocR8r9YM8CIDWnKmsv+AiltVpqFBc2m6WJTWy1ztlNdUGO5baSP73B12mJws0f8wmVQ/Y
kWgz6NMopwWiOvCeI/GXU8mMEFiv300z0+6D8T7JwRc/Nmc8skZKmGssUJ/T2d2yetwPdESDpZBx
LE+hiIKRTD9+oJTYmhoVRDfGUuKs/WKXof2Prh6ed8NfY393boD1tCx4gQDjJ+gwyEWljdQN495O
oc69iehKLOu6QlEpdTKTAkFDGOlGtbo+c4nY9FfO4aR1fOVcnCf2b4uERhY4gDvjkKM6+FQIEfCi
BkcDfAV/tre+AnOTXaSYcP3EHsU0CRPdrbjzG16RrzjIjzDNVQ3OlAxP7poQ3N4Jxl7tHafu/94x
5VsJef+63pUrsxZI6R1mEHaZyMPOWSKhcd03sTP6BCz9dUR7KkEw2Gv9I0ThqczKDkKGxps9PJ7l
hTqCs2eUQEHwpVMRZltCfeZM/UF7wlFxgQR+v308g4rbryOjrlFqa9OAPnIU4/o5RbsoKB+An2oI
Zunj03t1HGVGDptuh6yDEzR+3/rX5UizFihKd93fbTJUUJagSh/IOn+19K8wFxNvBDlHUrTjhirO
rNMgAUVvCnpMcWzSNHC4xDZtOVTeo08HGPv5/uL1/J16b0r6rl6TSb0t81/C8X7/kxTykC6ASIXp
U+XuzdlPMH/aSowC/2azwo/FJyRI3B3JmO7TIKojd4oDSeeGivk1jWjC/FTDcwm3E7vCJUgUYzTx
/AaSjQNHS7ljIqxhOxUGey8YhrFBW1jNCOsgW0ypZ2EUh2XU5oiP43Bkjp/rZWbzsDv/B75NgX/u
FnTj4hVqwDjbf8nYeOrInc1YQRQRKPfphq/3NOfP0fujmvERaulsQTY2e0sNHUyDpCPPmc1rn00S
mdjOTMrJ2ANUEMb5l1CP5/Eka9cwKtaOV/+o8CG8OZVtY+kgCLwJZo4eKn92uWbxeI2w8sMlAV/i
CkIFcTzXTj1skesYXS50e1ggTczJcIQrEN03U070MtoLvWe3nfdRG1I3eW1sVYntiaZeEV6/D6J8
9POlxQ5+45sFHp6+TV7jFXMqpnfHKUJ7ALvPau/6wpLSUsvhzRSdEsU0t1q/uq0+PIxgpjxYjRs+
h0GapgwCKmRl3cYWfdMz1nqiUCoRosoBSbPRNbKNDJ/6wmQTyjAfx8Uiq4hz3E34e4fQRZ2rDsre
qDjKKsbr41wvW1hRC6nnL7USeVyY0+GwBrpa5HiPxv55okEWuPHFINk++0RLZxafgnQlK1sJK6LT
aunXAI4RNd+c3vUcXAr3CSn+NjretbkdVCvNebsY7iCiNoikgkq59lo7BWKPwqGumQpt254GEWsr
RzE/G/bd/1OImpcP4wGh0Wyeu9QKJ/Cd04bxTwQ9ZXwy25A3g1OQ0Vpzg/lf1KS08CzXJsi8Cswc
kFjXToaeECzVkRIRPCiW0SVD1/Awi/3XfJ2RoIUDEX9jKrVW8YVsyYVA2vuZZygLhg9ZfF4jAMEW
xfi+l/Eh4o09xDmEpcd0bf0ytMh2quESAwc+wnkxBUErUWgMRgTM+iHyYbouxhcCQLhz34bN32F3
rpFEUo7RDV8d65ueVGn4O6lSCYYiiF3QzF/heimJRmvmmEF7oh2CXNS54NBJtjXzmGOzTS5strRn
V97dDUPILLV5pKjulbfNEBFRNEvh/GvfNRDV56/vvaCAcPQj/Nw+U5GgVJkJQ3NNyZvPdLwNjau4
ZINqGm3fiaCFh8tyA4VaN5eXJXwkN3YWZLI1dktvN2QpA95IAfXWeS/8U6j4TXlo9bW65xp7WfoV
tFKEpBaujxZ6jlMzgQ39WMe31oP29ctcq8WyivbV3vOvafZD4HRaRFUf03Jr6uU0v4ysFBONuqzM
78aGu/UiI/4BO/wgsrzxFxmFm8C0EohFovvsXkUcxDtllnVL+kDaQ7GtfWCgrYKChf5izGTQpOBM
bhCijDT8Alm0l2VMubOUN1E4uxoLzdOsWmAjmGAA/BbWTpkgcjgfTZf5MMjuYRSmnRu7U5XyaLDV
fhUqqAYdNo3/Ai4oHANo7/z/q3GT9rEk65vBVy07SIZONW6blx8KZgGQmGON7dWhE2ERYze2tCZy
qSRG7Vpsru6DNGCbkgnINh9zTeQWbFnjtdSn+igILkiQluQL2f42GUWzNt+tOVUPv3iVWlA4FW/a
RvoLLhDtlBklvgPEQ2KqhxAontaZO2CZvA4jN3NRKbtdoQbwFxQ4LHpimnQB2xHgrEuXkLjfXGGy
gJqt20wnLaKJK8eeiokyMkAN1xGXdf8pP1t41lJWr7pqfyG0mzlqbaogqiPXMN6/8Z62dWEf/uS/
AD9cIo8uMbxHP0nx5fk3jKZOMqzwoY3iojC7mcku8gqE4de4ZDA1NQWZs65Ycf/GMj6SfMc2hrlS
X1eFI+ZMjOcL74aMbMP2eULrG09mYPnrdiideelqf4O43QXqo0vi3HSJsHj1pgPIyzdWIdo0DeqS
cmve40hn51nyyIBURFcLu04jxbtwl5blP25cRJl/3jnOya3Y9j4LSrud3VJvpU7cb9dz9tiyhprk
KnCzuxCB3RlfE3k0wAJWi0gUyxK66E88k9BHmZv4ImKKrfRxX7AQGXbh8AGTuJtFbEsgQuioFXXR
pl3f4G6vHkJCfTzEPmDk5fzdMw6wVsQCS4A1tptogjaparI4eqconFZ+KU0D+nKHrNJMcAI7mOgC
HNrja76zSUjh5Blrtt/j8a2X2MFdAP0Cy6LcBTkatJhAFZzJ6pTKjjdAfVg6Ak4gqPtiEsS4vrg6
NRTxEWtkseCB0EZ0I/HCmq0j4u0PFmdrx6ynBFyfGTMu5uWiuLZTbQDTKBb1PwvmA25lkenBR7c8
8CAWYTFFggpdjTtf5VaL5CHXXeog800EP3kaewSo/G3xN/YIwA9BUghHmBMU4L/pST0lSFXDbP9c
EXsu9Uv5sK3fieqFIrvk8Cw0jGjNhOmbjG0jneH9Yza0AWR0yJCGBWsgsjSLqFVVNbY/oltOvbgU
xzgMiX+p1VDG+tucoBgV1KE8JuoQ4CvBfp9cWquASBr8ua5VthZYUdHg5xtbyI5E3NiF6dI7ryAK
8LIZspZRgs2GRdKPMQ8KS/cQsskRwUF1MnkJA1ysqypD9uLJazORE7IRtQVKsMusCrkbvk4CJC21
+Ee0d45sf2oXycpYxv8xuf4TM5jSlYoK1T9ySjAhqbajLO9i+oDvt14ODXUGig++4sR3qPUtew4C
peCfY+ZUembthHgrDFW9faFY2n1gYAJof2RRPtf1rZR7kdEkoN97gsgm74OwOvbKqm1bWsmJQ4Tz
s2+MCdBYXqGhjyKAXPQKdHerIPMOj3F4d9DO+6CzmRq7AEQ7hT4IBoTCQl72fRmxx3hz3sfLp0tj
dAZ9mUc1dTUphU8JSe9Hjig6GNGIchGT3/Q89H3Z7DkLxaWxPWoPygMEGRZinHCfob2tqJM73jRh
TXYbuYF0XtC0H45s+X2R+7rSUW+8sJaURmHgKrJscxxrlWfT5kBw06/Mnzx2CofIBfYLcTHmTZH4
tXpWvYi5ZzFolkuejqkc2T7JHQKN/6V7pLqeoF9cZxR2oa4i6+rVYPnm5CoCykLSJw1mkXLB0HVp
fLLbxM5VUoRUYGBkCILk50Oi0L2VprLeKiEoP0mpGlcJ8WGClieis4NR0A31KsLDnAq11MSzZaRE
VHowAjuuZLZcaPvo2zXfeQZq0y3WhHricdBvN2ClrY8VdFrZuP7YbwLSPW51+sd2m1V/4Nb8RBxa
AMK7Mi7NKqU+ZvCEGvULMbR9omICNnTOtmcpMTmGCoHxh/6hxW1IIZFL0BccU955uIumUQxUqE+L
U/O0+6WQg/43EAPRpwPs09oLpEUx1ClsTmlyeYwex4ts3hRalZ17a+7hgkxlkBPKGY9W555fMRDQ
QCsMuxnX7L5GXF296uPfSxRSCz+bOQqh6xl3bWyMVQkG6LevHzf9kiHm9A8UKZF9GfsEdktWz9cV
MHvJE6MM/bVm6rLM9xnZXRN8MTD45d2CKdENSMUtuecPwkxg2/KbQtFYJVkWZ3Qb1f5MopIotcYM
FygJSkMWF3IOtB6aQm/6nX/f8gUZkjrdHDSrPWH+eTclGkKS6Yapxni9zjOrnfSpjMmhYfdAtmEM
G3fCTm2Yom71oGfVspTTCOJdaSCeTSc/0ChMUQmRpMb6kXqy/knWoVcWrwTMS1QgzuM51CwPhcsJ
hIrWIY2CponJq1y/RL0N3sWvTnzzbuQsmvDivWdu2g07ofVMIt1XcFEU9cDdhYOF4MEYzFNzqCgx
mmF+Rh1s90KuItBcfPOej7ihkVLcYytbLquZ4jiseyRTeYeFlf+kBK7vGIpd1IG4vDKjSWASfYXM
DpFvSDgx2ZRoLLRJ6nOoe4idKOQ4gwpD62yEIv163CB0jGitT7YwFVqnqCImpXtvDH8ZVT/IH1E5
A/7JH9o9dpHXarpwNI/C45r08j5ksvArDO5cghEak0CL4GYQsExJoPGVcudx3Ywcfz8hCu+bAcOT
6BuuWF85CQGox9GVEz0BwGmt2Ni0Zp37xFaC+PNjMX/ZNDHh0lRxcoaB6HgCMd/01wovmwhsE6NJ
6PS0dVtl8axNazLaQTom8J5YqLVoNEU8fIAiMHhDyvtzaZMmWG8cQHTEG029TTZMyKDNiR/rle3b
cJNJpRl3uIXCKKQNiIl9EypQix/0IYFwGHGS8LGWLgHYc2kUfrT3WkzzxhthLbyi7OesNSRmlf33
uEWDAx2Qr6wLBlXSnKx6YxC/b+mAQlDvuFqRpkp2KfGwTmLthYyJ3O+Oh3xN+YXcbB8Li84q2nrU
o/WvfxzBXoq3ce97op12chNNxhiDnr4UrtTiisc0SBc2jlTyAqXZDllqwLfYgAtgIKomDffqF3dg
2pF6ONzBXNeAo9fxXbyfe/8J81UsZjsUOoNjVkbg1tYrsclJgYDwDGpBiqzYTid+nb29IvdKYnG3
yF+Gu1QQlxHnVOhziw0aHNSlWn9fN7YMIaTuJOZ1EDcUNaopGM4PML819MvonOZVGb0yzygIHYcO
VbsBJv7EBQjcjX0UJDNSnlbh+wcd1Z10TP47Ee2iFObB5YG+OYlBrxacBPMid5HPP/g5zqfZ7IDB
Gms+GTsLrTwIFPCuEMWS2JUhnucc1hWa6UoSLXec1Xm65IWH0/mVl6LhtxKEHf6bhIw7RMB4ION+
G0sLfrErjIJTVc4ARfeEmSsAokX5kg/nFxH1cZtqgguioT3LgdPOhEQV2qlt+mzHFeEo6eTd3VmL
XX+ETvR/O9A4ozvUJaOymQOczX26qPdsdww4czOSNNzclG0+G9UvNHy5mvbPgyhKKn38j6xiUWdk
kyjuCYR6IpB04IqcZK8ybdsZii5PRemmx/h1E1jXcHre+EFZCjdwonmjxf9UfXRjXt/4fYhWU/nZ
xezHAeyAFQEGkZu2FLnB1x4pA2ixgNh8jnPhyGT8z9yWls+4Q2u9RyZ5We4fwJKXarg17p3MID5R
A1adY7nyCWm7T/s/gV3iUyi66fHGR9ZiRFi+7goSxlGbR+JOq0hpMbFh5f5nEQoG5yGYAvb7yF7M
Q5Oy1h4jbfVFTIMY0N2WRHuu7+rXexDqN9lfZhFLfYGzYQgTUqsSLPd3F5tQ4xsa5cnsuu0H+oIp
oWS7XHL8cScrtsPWkQAW3zNM0PoyCdkpk6HZdt/SqaggK0DycbSfrtwU0rkSB7s4OI7UfUk4Vn20
tCPoq8tdE8zfyIl+1PwuMpIRwc8/00CfloVjshC+9gmebBkAaxB+3ZjZ3bp2NT8PWbeF/Sg5BQ9e
pHBWA1YAc4Q8Wh1/EYDz0zzIl9vq5BviSLddF1o0dyr1YShjcrY/VZMDe3bVKb4ZUhVvW+gwSAOr
zHlQgPz4XOQt/4Qy1X2N61q+eyh113sbwjxmeIFUke535oemEoIXw9wi7KEnnZAbUS8OYQ6xBGq0
6kSUqftIGAVf4alFFTznC5jKnVrSx6J4xswJQKFeUOxgKE3hDsTyr5rl3+qf91hlCfEULFF4ayHs
ih1SVLV4QLfwS9eb0QLtX9uwN16/hXnKQxkiHwjLf2I2CQLuotOp3m1hnXN8nNowWBnJo0j86ajG
2ztvAaMw3t/2bRLyINVxmmRe4AqLhWcFfY3PRLoDcNzM8MtOKp9fbbAfXekuUAgNydoeSpLza8r1
2iybvMOI7AsGqvEgXUJlEGvjGar/hG7x54eiVvHLpjbAS4iKzBsDwFLfFjw/JS4r8ivgMbvIBLEi
cfSDydAh3lRffE1q+LRNytSX23KX+JJKclA7Bhxl4nbj7I4Dq5gZPQ6BwfH8gxlswhIDWRhqxjwG
g0nwjPc9062H7F63/8DQZ5VpafSXnrnkxDi2//mTssmqJTT0IRNsvGTqr/GNRuN/SblLipcUtzRa
UmbZuSCVV/9TffYZwfhMB4kEcHGKdCMaxWTqkQYCA+U+f6rblsmfpBuBAcVgHCIgd1mQ9DrsVyyx
K/GbAA1wgqDZERp7X1H6BiuJXJYf8BUnVuq8xa1UPy9Ww2bHYosa5Y8ExX87yXzCPEBjNdtRVUfc
hougG5ecFx1FZXsDU7LPi10rx+wlH8NCIe0c1V+tymWiwXshFzOi/UuJLdgTycfAMZsnnTc/nZrK
lb0nEmcQR7lnofnP1JeLuvT98/DLGC6w4sOeRKunKeTIbq7siSTEeD9VKlVRPQsSTwT8EVvoHgOM
LGVOT4obWsf2Ncp6OvW1aroImSMzJGJtuu0E98BQteDbVflIkxcNUgIEc3OibPzdE4gBBANqL9L4
m4wX7UsP3DdopQCnP1z7AxXPMdP9e+6EmvMktuTTg9+CsrEvH9aZGduMsxmf8Zwak+6y7Y95xRxY
X+6tFVnbEG55+SU82qgUPyfzT9JJZEycuKiyLvQfor2bnweVVgFaJ/9fFs7bcqmElTLvadNxImKW
X4xauPRQ0Q5Yc60EYjF9FXWCKBHOxQgIo9XeoXvNGt6MTisHfAOI7K2E/30GDeAOu4JNGEYw7LMN
dp5dkZgT/1jJhsdeK16QSez7IS5c8Rry+MBZMJg3F9uabM0+IwzP/rAsA+2Vvtq5gbr9bo1oOqdh
Vbimd9tntO6hdwh7ShsqQ3lZLqNe0iMrCrGyRf+HXdkZWaRiA9a+t87hdBL+91gCHtQuNPNP6E0C
b7ubp2C50wF00k+hKBzOc5T2OE+RceSNd+nYLwcHVhJdcm+0HHouEteUe+kIcd/SK0QD+VThOw2f
85FUHoOBH0q1GHx0MQhHT9fPMn0E11zoWyf5Yvxsa5yJMaFjXEq++2rSb/D0W33tB/z8fZ6ak1ql
I0AjLbef+wNn4f0c9HPAlESRmvRTe9sfb7g4yDgy2Tc7LhG2MBeWuN+CZ5G/Ht7f8L/8XHhkCazu
RF4QKawEaEpEUpKG1rjR2U1EbhLPi4zF5UdSg309VyqBeQmLXzwhMKYP1DjiXiCv3PmCMD5uy7dw
8WF15dPuN/XLWw1Gj/p5ORboQD2ff6baNvK3lSFRwP5DD74qJGdoIwr8RZRF3faWRpIVDn9wok8u
OXnjhYw9TAbgpcU47Rpsxz+ar6eL3zQ8RlcQ13HtVMFj7ROWPl4Nsq88Cov0bvQM2UBff385vP9u
Zyz5FA4lB7Iw7NSPJCAv0GQfAJ7da44nGGUCBRATgVMvJSG/mSR+x5t1wlIGw9Iok+MGIty/Tey8
5FjMF5NJbtvbpaRZDj+ZZVUimAC+iF5S6JaalO3Kbzx4ASHDA09CMBdQ/60NnCsYtf1EeULGflYF
KcmKFmDqqWnc0CirmQR/eEzIIhcGouG2gkF6BfcrGOh5J4tiYmLLmxCNY96C+P5SSYNOB5TQGK3Y
BAIfZv+tug3x6++2HtQNV6/LWMakLkI08SPhz5kRLNIG4VH/mgKU7OuhFZKbFXcm+Ax55qmeciue
86w8nrgma59+InAUat7IdDRlVwpH3g0lRcbFSuIbPDM9n5PxGXCwaEHr3XULq6zwSI68pgAr3TvH
CK2XA+GPk8yes1lmA3/D/yQ7qdJMV0/tbjAxhMlCH/0DGeQGOJq6OIb8rRW1Fvilmtc1zBd6TxOs
urwS41jnDJRFY0ruW0HZaM6fBTfmtUXD+h8/5uOB1HyCa5lu83b1+lmupaX/gUBJKc1sIiWMc1nd
4ma8C1tO7jrfzA6M71Ru33zbzHANVp04qfU91Fo2+40cIN3KSWLGbRSNGp5xKmifYvTsawUTrdDK
nYsAL5ILBZe9C0AhPv6xyHJl6xv1nqbYG6r0ZGRAN+5u2xEMnaHaXK9Qo+kmxCVUaEB/8N7UB4fL
w0QmiF5sJOI1/85Kh8lA/8gYtMQ3w2Vr0iAaDwuJa7wg9mIREWyx+EHJ6PjYKpVy1TxwGhDuKF8V
3oe8RzMi4GJzNpCABAGGOnA57zWPjCCya8FShHvMt6iphuI8QqCsRzpQfbASiWtN8UUdHZksj4Mj
YVCeUjktvTrBVwywC+UjxeSYD95txIXRZwlJDUl7CbB0ukSbBok8cNw2wgCpot3D0qo5MHSgs8AQ
3V7gh+g/XLu3/bWpuYCxYtEbymjwy4KCiSO9ohX/NFNFcCcWZDUmOd+MSPCd5xW9KV4Nmwj6vdkg
dW9zZLnBTrtzBdUztS1+Ng67WGK0uBMwwmXwqLpOaIlmR1vlSZxNUEQnEmZTnk53QMLtVXCQp3x4
wmtnFlW6oH2rmQvlInlqIYdpKKPOfUXXqpo+q7c4BcwcY7jPKdrc/hHyvhuVocUHSIswyAkr+L04
3PsK0k0IbCDwz3TCLHx9EnOnV4OGdlMsMbpecTe1lSYaDXcDQYKJXRE90uXY8kXO00CCKyf04fUJ
X1PlOlbFWaZcREBdZuydP+XqBeXKe/PODgmo/Hzlb3QkEpFSFCQ3x6TP5u0DorKZv873hMOMkDKg
GcrcNlDMZ9Ge8NGI09zdWiNppPxqOJvd6akC5v+Yr7tdNSpzVhK/Wa7aCeva39NZSNJfv6xMKcPI
C/SseS0m9G47usDt45/wLgQ0mGbhoIvdCFu4Ps6tKCHvIJTlTAt00MO0lhTaSuTX3ZNYJ5+y0zSS
Ivh67GyB03CiWHWWCkOHZqDRFj95Oyg+CNZuz6kDn+mR5NWssbeHXdvttCAt3nsuEglMtFdGbaxK
Z8ls/V2qm8N+CSzv1Z+II2KVvwcRPKe9Ztl5L6KAj4fvK18Md/jmf/nOz1v/aCi5a4WSXVvtttpL
JSSEfo53H7eYx/Uv6pUZ8JUq8cB0HoeMTDcjfLTiBQHiUofslZ+9TZT8cyYxTDiVlm9anhmx/4Zf
sPG0aXh5sGbZYqbB782SARJV60QYMKmUVjAVNqQFc/MXY5baDHqVNEmlpMs8GZ9CmceCvAP/UD2Q
dFUKNQ94FRcsjjt1L9tTtBiWdl1g2iGjLoaFUSdB1EFJL95wqD52QpvUaZhCXUtcKGkEfTYR8cOF
RcctiGbHY/dJFqfJjb8hfK5yfoop4kKZAI/h2hDj3BHLMQn0aIyCnLM2Yn/EUPRIODQ9n0viYl6K
ZbXq012WLWHNiiWO3y1rpOV61sexDQVmGlR0ufN728KDhH5JS7E5MdH0J7K9SDFTXvqHjsKGAaM0
d4lJAUhd3eMrjzd1bf6tjoZU9XfOINwuhxS7dPGe/6tMfbr958ThDFxtFx93EaNda7NCvmqGe8es
Gb64AG0YMFCecJFhnZw/AWeS+0Ii0yyY/Ky1vehGfxmvF+slWznY1QSGw1nAOsCAeb7m7K2aSovc
E0wCnF1zNszkhs1V3SfXR3Q4zhSqOeMnjtoB/jD2l7gjKS4+NOu3rkPn6WlaL/bJuZ9t4ZR2VBqO
enrLlP1d9o+73QUGY2Vy4q0UntK5SnrMFOJMEIw2ZRaERTvBm/Ql2Z6wywKDX7PbLupgrieyhcfR
qk0jJuT3s8uk8uF9pY3XZuGkwArZu0e11PmrntcTW2NXH2kdfK96ch7kAMfyy1ubL4fzmpdtgL2o
a+FpsRomPu3ZLXBkZYg0sr4ZXE+0ObSM3awiJeQT/FDp7Yjoi24stAEWZrEAbaplO2L2q0NN9v2r
An8ZlBtlczLJl9p/ZEXuDpaAJ+2nrdhE9SyzVbkCuxSFHychkSHwPba/oI7Db/of6TepipwHRzOZ
ejJfUPezlDjngSsBlrvNtYdX3u9HCxIOyOg3hEzgeX+STDrKZeOaJk+lJwTkZ/Z8y+k4nuKzXSp5
vx4YIJYVxg5NoJ9x9JDz1ZNSpGs1I8lCnB2gcUdnF3FnsgLDljghU/x0UHeZyyK/Y2LVrl0EDNbK
u1u8+DtvlPa3Ucx/SJ/pTP2FZv/c5NBTr2cCGshDCpne15TofPIB1UFPqDmaIQ7gB9UJ7obNrUFX
WT0EEWEK+tDygTNmGdXg6fGqV0gNMjnIt0oRWEtHplVBYrpdXwFSPb7XnL1HAolM1YD5yjSjy8+K
itpGkTjhfG89xdwcvnupatzV2CwkwSfS9iAtI0ID9bVTMB+0sqG8zC8YrJkagcVJ6PuXV/RyhCV/
KomxDJVs7JRXuE4NAexGtgrjf2BGZcm3L22GMybzfhRyKgNx66p7go9dIHfoDbqSWf08o69bKJS1
s5EKicwV+PXfM53JGYQzZzhNw+tYlhR5PJ6zuhx6n9uEKipf2YTLMui+C+Yw7Iu7VqBig0w/7cPA
0WN6bVr4eWxqWLEosN4VqfN/McxTIjYDahfZN0yuJr+cPY89WL7ME2Sscr/7jf2U3VwrHqYHrU2H
xNvikDT8r6y3FaoXSHIAf5NltbbenUKv+3OQL7fuxYEDnIzl47wHi0fDfaZp5IGUcZnMzwxQ/Rez
pN21OQmdGEwOAJprWEUWOSZn0JL40XyKhN2r6fk/+3IFkY65yz4ql0Pti/wg/t5mGoxJ1TJBouEF
WPdJ0jkDFPPU+FdsO9ixJg5WcYnCE5U7HjST4bBW+odhPkagdwiJ429897tjAwfpWJjJmiTDDPbR
XzpAU6buR7+QGGc9Xe/hAPeHLN+SoQAbNrKVBP+AhrJE0ldm6Eso5St7xsz+uILx33WMwiuuxqHd
g9Cr/loWjah+H1YZu+4v/2Y0bSIMxjopigwIB/vM7W4WOsQ9jJSExx0x333oOUPFu5v3YyfiBTCm
7RJR6YwEG3SvygkrgiLjtg/HYD2vd9G+j7yneyEnCvkspIT1TfzcrOp/JXPJaiv53bd6fQn5zFzi
3JpdZpfTIgsL5bj1t+akd6a9yHmeMPeqH8sBQB2DwO7dqoq+FGe0I4iaGN547o8gHDnc9XP475xo
Aqr5z5Bgs9XLLstufRgBjPHl6CMuzsSklFFOevl7mmuOhfPAnXEyAwS65+3iD1X1FGlIS0GcnK+Z
YQ2ggGKMWIu1WbsjaR4gTlGgc9sBbpl5Il3JDHTJdbZPTI/jdqQMFaxQtjWUdDPSzCm5BMfbJtf9
/0x0E7iF0EViIPNMb8jR9pVXCmqyJJCDMmVp3+z8IL9yHsld2Vju3du7ZhRaMtWxbVlmcVJCL+lg
faduA1Ib3hqghjIkKgUaiTnrl0xVfMKdD1RPF5ky7ON5PIEHxXb3ULsdTYkCxYlpMgO9usFE5atk
BOTNHGv+iChpc9Pp6UR0bhg7pBynkIgVGFjrD1RFC0mZMswyP8Msw6chWhnNVny65P0z8WAtFPkn
yvcVHxyN41Lw1ulweOJcqSRxZ3swjUFFelRA9Y4nJ/1eph5LcU3/qTk0Ik7Ywq5caNbv7njElcpb
G9EbzqFBCU06dntVcAEf13OgTL6QheeT5UnaDsLFTm4hN8lsovcYZwu59lxkQ5FHfqqJdEaEW0st
hI6eZWieU3QTrOpj2HwJYx8/VGnvMf/lyFkibNCuzxeqrvTXq/C12QL3n13DuAy5Tetjlm4eUmkN
I/HQFDS2o9EqzDurBSyPQViYQrl/1nTwd7DQzIfFyHEITtk6zTq3d9fAR5HPcmeAGtS3xiCZbjgq
vqLqKdpfv/itKmWYY2FqRyXrOFeZAgU1naBBqxD/H3uZgpCSP3hXdDn0gqW05sK+TIy+XNepYVbS
tSkNXu/GuqNJzd4dFKZ6SxhbHQ8VlqYigJ80zWp4YmhguwkaAWwXQe4z+WJ1L2wCE3yXNmPuFRmN
g82xhd2F1EV0/51sFiT/2olEDbHnYjtoWHJx3xRIp+h2LdI3zXTxZjJ68nWCLrlbN546+W136Ygd
wFY0szEg2OWTzsEWeuUl/SbYlR6MZpbJJSy4orERZLi5elDOaTgVa+VoZ+VRdXO2mwJrthsFEv2d
mvWn8h9aauQHUlfLiUWwR1acPo43h6Np+Oee3IgQGyWMsueqpdE53a5LBOqBFseyn7OUlpo91OXi
rFYa4Em6KLO0RRfWFj+VRU53AQ9WlHG4gWp3bPhuxy607vhYJM29IIA+xjTgEbcHIOvc6cSJiCaw
DCvEa8k/2yPA9SeeFF6IOxs7iX9PyZWhCtXhrQx8siYxQOcpRy0Cx8ymbI/75vCVg0X0JWH5lpeA
r5YhJXu+ykaQGfALGyuDHeWBS7dOsG2AT/g6pimxWOLVe+x+M4Ca1anRrZgs5e0Mz5ORwVYLnDU2
M/Su5c8v6d1oJrTcoyh3Kes/tLJh2ni8OIgetAngrcRC+jWN9Xr3rSh14R0H2diRi8wIwTWbP3MW
39FWppxUGB/ay4wTbiLMJoSW20qZb2wl3WOpbtGWMkVZJA19YHlix4yxU9K2nicoirYuEg1Xjcgs
jA7HTZbpat/4wJJnNa4XtEvuFzQeGRZFjyIEpvSSXEkVZYTk8ACt0rflcU7EE1LYHt9k1D0gwJ6K
NfEW5McEeS+YSfnQET7IW5QFLMm1PKDQzX4yaemo9Th9DOI3ynb9ny97R5k5zdDq0ZTGSQWEKXt4
L+ZdqwvQSjyYjUr9cZvoakKVCR9zRTO/IRHKJ3huFNJGuV9/OJ+Y7iOf6nWATLEspPsHcIUeCinm
QxKPO68pFQzat9ktF6pi3AnRaGd0yjGuYwMXHg7kz/dBsQ71onKVeGChZgtbEVZYrOijH2j0kM2x
D30Qk+mYW0rjo/qz6X8Yvcpr+lBRsjWwFXFmpHfbKNaArmahHzSYB8lQJv/a7LG2qm+oopdLxlUt
f8VA5DXQNwVVPctjTicby6/TaTjkdOwTWDgW1BpyPw7GcbrQNihWS80kAlfwKof9ovia8cjr41UK
nNPm8kKdgCLOYQotDiYyD4+GMajjd/xv7oMtTaFQizDRvwI1XGuGRaGobsZGnkk7tvnaZufwdPDc
c06JDYEP6/cmY+nLdlvCZE6nBLZ3qvoCHuWevO3++z9olyXXMIwcrSDnbNfz+dqX9CmeMZF6FiAk
JFHoe3TzlPlShGeEU31Lz4PyrwX8lZ5ashGXhROvQkkYMgyFLjxqLoyBf4q3pG/z6PKYm9+cLZHK
72pmJhLgph8rp5ujwZBrQY6ay/XAWBWwcpg8Dlc02ZrZe+M9h+AphZjt1KODxLAIEDZSsnSeT4LL
m4C0YwFqVHRLCpnVpPWX+Ynrg0QqrCv4ZCPDVEW3kOc6YmDei+4v1B3kWjlhgdxrvaNScEHX5DBy
o+ILqvvErWTepSGRzgv3+vvukW2YWBhQvh8/MsCgHRhykR5MoP9yy3gNXJBLqD5f8FOB/cF+fK8/
+uTuajYxs8xOfndZjmQZhS41BkzVfni93zrzLWlLBi3MnhKIxfg5YQp7vJgtqjdO3XFhOt5W4fc1
QnbKc0BqDep3aMeVS92zoqTBjVmqXwGpZ4roUIG/Z15hUrzzeUCVlDRQCNt08Aa3wK+94sB8ySAK
d0qU2NhbzsExiRi1XWVt/AX2BfdPJHUwXJjvVdHMoH5cZiW04ANspac91cFdSDFlSVaTlWKR0gpH
QHTtNDGtrkdrlE9Log0mrdn7BHikt2aPii3mzreoOnlKs8m6epw3OI7ZK+SmQSlUSfhK1XuLbYL/
2pa8WPtWmAz+Bu8E5VOk3NC9LyzRpFrybxx6N6NSi3XfYBi3CEw3aerIVDQ2VN/JrLqc10gS5bmZ
95peE2EyBDgRipX3eeLIO+xcbGNuSPqRgdzMA5dcL3o+x7npMsc/elFiB2GhRGcm3q0exI2WbUns
sjcj7NVZiXcIM3hBGW667EP9oS8QTMToHaamQq0nxtgfUc6yDW6ql4VBkJXm+jT0KdiJaOR/BhlH
WA33GTuG13otlkyk9fTCfkzd59uD+iDOqZ5YvWm/hauQg6oKL0P+OeNGr6Twkvfbfacc0IFh5iZg
LDMBtmhVFuEALP/662erDAv/ngGdmSC99c8ilkIrpmPWblp0SE8nLIf1rJ1ltWXYHUgaW8JRn4Ii
NUDowjFCyRdj9EtAbdpQUijomd7HUa5HgwAK11nP7wuL0ij8ouJrVsDTdmRESiXzvCFGmw8TNkGO
ZAm8bLh6Ku+ZB5bgUJN7aWIrtbCRlmxmp6MM5y8ZTGnbTR0Pd7GPTVZHaWALnRUab3OcF62GtWm+
CxsNvRcYf5qUPzRj3Tl20bH0cNg3RSBJjgpq4UeQw49DZcwfYmMAQYEH6O0J3kMwO/Q/SAODvZUJ
HdXp2Kud9OtbzIrD7WIpuiCm+bVoAQXTcUH/WDACsKd2QiAcAZ9lyspMyOi1ns6j8TQMJNAcVE3m
YnZCZ2RdpjFZ2HBmsFM8Z7oki001uJVPO1Z+NvXtwo0BEqZTeIDvLwEIMTftan1WIILAc6xAdPhI
U3iv58UlLUbkNKF5vJqNu0/x2jwiYWkRXL13UyUA7xr6AR+rqr+nklpGYcD5JqNhTiC1skb2zmru
6DKNWCAKQ0SpCh/rWffDWCGOby9Qr/89dax8bXiS91od01629bxZbeRYF+gyu3KtZpH5fW35AN6b
8QjQbyByataLSuw+ITPtrH1YtIGP9X7ijR9MOlIkoamtu8uqUKXgFWmU9mxDpD4mkPGvwceDi1ft
PG22rszpauuG4q7AZNdtx1k2vW53B6hXN39GU+ZRoY5k4GizBns5EGzrbbMqtpJXoxIVRoAB+Sb+
ArCU/O8YMM1m/ZIf/7MUBPOJnOtGJztTHS5P9kFdAOZZvqVe/WoGMoS3y/J3hGQe32oDD3HW+Oy+
xbA5M2Koq+CEigPJfktDEAw5daGvUbhE+7ueWYslEzKkrBUJG4U5VRU97vMVzArY3F+uBSClzcuf
/lRpoT8HfCEP0Y4yPvrrn01ncgaxOmtHeVvbx64M+lN77EIQppF8O9kGbliXbVUPX4fkkqgRK5jy
X+pE3+pMMvsU9dhAiigmXWkO5H94+vx7Y0AJ2ddOq6Wll7ivc059KVWMA05g58Nsm7p9ob5XhCKl
uayxZJwKJIzsSeN0sFkXxFbSvPwf2kimmayMJqEp7BPQ85/CiwylZaAXyL4xnBZlNn+d030adfCl
Zh9AGnRBy3GQ3P76mEHjaXbDg3wAdWsdJUpOJXPund3eZWf3bUhWhRbF14r4HmW69G34Jf6FkUpn
F49Ns6lXfyinA9I1uQI1QxkOsh2R2BYbJqn2xpwHZe/JZdM7mbWInppGJTZnv4QRaRfp5oOVT5/0
1XNB383dxiB2pf8UJ5qPJkf8yH1+kgSe7loZ8PK1seCpeQpsp09V+EasCWJJKomyr9PypkKxDihI
ngBzJ1mpGrMt64VSC5T7ch5LOhxxv4kwFEVyU4Z3ETM9MxQ9VylaV2t0rKlBDKx8iybFxi32++Ed
7emA27S17SuSFgedeiv5N0sp+Kcg/Y9nk0fn3+stSakf0nY5Bj+qqVMqA5uiRGZeK672/uMxM2wu
hAwubGclnzVL0G3xyoHp/xO13L7RU6hL6gVu0Pu+uu4oLB19mXzpTnwTGomCve7Ydro8Avxo0YHY
TsDzs4XAjWtOHKooINh0dtgD4oG2GvvzjLuu8QOkDidwEqwqVFhSUuYA3tb+hPwiZrCYUcxC6BzI
gsrZ+9GDlrPmqt9x2vYhzJirAmLS0zGvk7wEE7RhXFRNei17uV0E5ugprW1P0fMST/l69/4G32wW
uXngx/cR/ZatHYnjuZNG//2pyyqaHdUY+eZyTWa6Lb3Ce84miJGSlowPJzv+yaVZ773DAaN94zcg
OeKranem1CWP9VuGBN3LB4SKvfcMrWWc2iK9E4P51i1ANL24ayg/TfqVJYPwoIp0PO2hx7x4ls5l
Er60jkFQ/zLwMp/VXr1CrQQOKKSZ351YWfYxZvwgJiB+8/1Rz41zRtpXa5keaNZpR6xH8Prx84LW
UAV7geSz6HbWS1z4igcN+a2fWS5UC9V/SZqT4LCJ05MKnQID83KdcDPHSNmXyriexJ029evu9D/x
JKpjAoSP1Zmde4cTGXlPcquMLCTCjrXfgP2ATbUfr7sSwTkX4WNpNm1NY3eIeENWNX28ZcCIIeJ+
sBr3MKj9lvP+9LJSvCsLxfYizs8dCZ38ZsjUpDUubvpX1cHf9DUZmf+NAKjpuL9cCAfx3BemPycC
YMp+HJcLOF9zSETXOxeKCHcxlfRPQqiYgcGjj6HBg0sbIHkbm+I8h69f7MHRnLcYapvuMGonigqT
f9SLrN75iB6CnkVHybvJy9qrm8Sx0mx9GNirYu5j2Y7xzRthr1yrdRBWDUcUU9t2IbiZ/5l+bod6
lddWwzVGCRQOAPPI7e1RgBgOjYyfTcOq201dGd+rxnNQmZDTbLC4ozVbeQAgIMr8bMOYRYr9a7FQ
gE4/o1iSJSU1VoyswwNHiMyTWF1frT3CfrkhxwqrmaaonI7sP2Vlno/tGRlluiHMYoP60M7dKo41
HG0Wn4VDG6RKxzhblLYYyBpwlkx1E/fIepJHx/y/qKRN8Cww2uomygBiKYIJ+kYWLmVxCPRhSHjG
bTnPwej+wTJaTszmrPb9dv94i0+ImytCbXb2qKA0wByg3+2IcBCMWzAwlb00ITinV/hmYmcNFJ9x
y0/VoGdX7t2n91bj6Rrxe83/NMZ4GVmwNEnQaD2RuyvkRAshW9d3AvdbfqFrH6SXl2JRBRcMX2aD
Yyrzt5fYzEvcQfX0ycVrJcjIHIacMz7wuhkIF7nN+PL/BPtD9qFvF9SeZOmZDNYOnbZ2Hw92IAh1
jMbB2uwYKdxIlckia6fgzNuPDtZ7l5KxsldaqMFQtdOr+Bvx07uyo6F9Nzc7Wv7aK+lBHNvbg+ic
9gAixXpk4EgJl+5noKaw9JSY9+QTqM1LXNFbsqURg3mdy533cVWezo94QfpQw7kWH5kvVXvGCMJT
VO0nv49tFBjEurgUUxUKrjyMdSIgaBCYcsuHYM6dURf6Xx9E8XBRQ+KkvPGtY5mVdv678/Nmturd
zrBpkMsK55ZnoA9NJzz4+bQ4bLZnlbd3Z8lIqr1g9xRFqt2KKt1xj4aoFeu0X8byrAs32A6eX5pt
jXvDYzi8SSPFxNhdOO4JM//+clKjF4Ncs9rILcDKciKMbZ4xg3BNY3ZvMy0UEeozlRLF08ou+bId
wY4cmBYXffMDd3bma0kPT1vOXVdmHKpuhvJ5r/AbQmJPFq6yBcHJ7gIyQQJgWToUx75MN16W440w
MigQp9bS/umKgL2rLW/lvlnrvMZ/kuWTBg+n6S26xGUJczecsAKQNvD6ujL2wBkN+YHcmP2UIEKb
4bOTG8LLyZT8uR6jTEWdnEwvsBmzt7OIVez15wYWW3AAF/i7COMP8TSgfOU+bU9Xy6V/rC/oF9Mk
5ag2XPZGl4EzIyVuirTgm7ebxQ2ZpjkT8jZMLnwds07RxhUkDwn782J6Tj2654J3l801WfDV3LId
IB2adT0ZbnursgnoKMeS1rBOIy4DFrLV1LTTqsvXTazM0kdDSd/caIRw+JbSl3eMXHgS523BSMZE
9BjqsDz85rXcHtWQ/b/mxyhzbjaSVzhY5YYBFib9AkLRDdJrJJAy3K5+Bn2JnMuFT1C/wARQzNV7
1usfwCvDppCovPsrh9TM0d3Dte2La4ZjU3zYCaZKT0bwvRNl1FGCBn9JaM542iks/0mfeIbLsWme
ac6+K+JXlF6SSJJmjrUoQ3MikcERYUttL5Mxtc9j8PjGmbQPY9EQPAGAJLebDGrgJoeHJ5qWGfw+
Y5lXRITJSJjWGu9Z2FAaXSah1G85zHdVATA7+8DLe+tRxxBpJi7oIZGsDPD1NI6YK+eh6ngCBYEH
Yg4vmtjzc+LNuqfzo+1raUzRJ9T7PKlDt+w9eOpxC8BAK/oqkXDpSTLsWChp8fSh0cdY6vNzqGaZ
GVKN5JI6aqMmIomYEMgPFOu0OHV/YzoXykqh0MGF9q0OGRoHIL+Y33d/zd7MiusaNafIiLWdAhKx
6W4WAUXGLMGgyVCzQZHXVuLIai1JciFBgW4YVOPjUqdZP5me0/c6LUJJCFiPapTDsGmk9DGNd6f1
PVHb4mPOh28ViyZ6RTrAdRrsCgE0GSLpv9khdv+/6ND4OGNUQFDT+b50Sqd4GC9eOM5LdFB2pNhn
/SXIgYOmQeks+dkWtzdgng2UPN0VwCPwQz2rKLQNUflk/DfsENGy0NDzopbo2w7nQt335sDtllq7
dHP1epiBtHq3f73H9ksn7B7akUcxMdQXN6Wy8y8wCOOinDkZGheFlX3EmKehznf6D9dqEMfQRDgg
fSnuhK7CT0Xm1cTRLVEtf0KL/OjEn3IWwBjaKgRiqrIeO6T/C5mxprtfZhWSZkZnAfQttmyNe4K4
RPU0amDHAnkzS0Ik8wd+GNfzLbYKT2KxHq98ezSGN7fiKYJ2lrjx5vJ5Dm8ZpxSOxkJaDYMN4Enx
pDvQjnpURE9Y1aIDGDFDkmPdNoKc0YAO7deJRIqMidE6S8vEdoPbmumgJQTqm6EIu1w/AmtdSZEt
Qhubq4hnCwB3YLbwhhEgM13xyuY8rMOhwO4mgxm4HxT+zVKnh+z5iVNKNFhH0Fs/aDxwZBBR3XZN
6V6C4uzeTXcq8de7LSa7l7YQ+a26Qy+ZESUjVhVY3pLH00P+CsAdptYWnTYBj4/zGG6S+50ncoUh
jNZu7qF23Z77GhE9eWBZx3Fi9lGk3RWRoT3rv6bU5HDt1sNniQS65248o4wek9bOHiOLINxLUS/U
eXbF41U0yFAbA/bNMGRov+ChYOllJpyvgaaH5pOb/j5RVklc9TGwzYG4stkt7D65KyXKAb6as9UH
Nx1Q4/Hv3YmT8onIqTGaFYBmJkJJValt09FOX5zFeYU8N29rBHt9asyx/Y6zM4SlwKlx3Uc9y9Go
HWvGkZCKNcq/LlasdTOfvLgQ6dBGdzjgcSUgRUnf7Wtf2IfEuYHnHjanjlSDr6ge3GK3ACiPkhdL
Z2SOImX75FqBP2LopLbEgpOjEsXendmtw5EOQ68/HTwozoPu0aU+kswS81qpwyVw0WUgZjdIpm7D
++ns3Y+1sIv7NTAiAEzJr4ZkXIeE3HghO3MhHgtiGaB0Px4fkqP3ic95Pl7++ZjOzUOdKeu+ig+3
tapYU6+/Cd+Zx3g6q2kxMmOdH1lVWM4JT5UvZ3aZvgD569RLyQA1pY9Arq154c6grD84ffniETHD
5cC7LqOvxmPh23CPIZnFOf2r0MstIsdt17oEH0RWhgFoJop2cvWz7FeE3DsbiNKbi3MZeP4a3Rru
oaCAN5JwTpDV3OJSiyGFi5s7LicFEfHKUvxYwKH9ZjCzd3AttdbjyNZO+VunwBuMgB4mh6m06GxX
lLjBl67iBhMVNAka73AznV0zpOxD229bXfvq2LuETdAId4VXK6qvrRYNbN17TrUm/8cNvLLCZnbx
5oAWkYHZypXp+aQkz63bjDItfNNYuYDbK6LCSty4IWUIwvcmqOGdTqB70GuS913uN0/T9PVFHd2F
ciGfKmpnZZ4R1S4jE3nc+yBjmw+CKmJZhCkWWEl70YDgHkAtPCdHqb+eOEsOP5vRhM2ky2PuJCrq
Bl2mxt0MX0s8m9jNOTASEFP//Q8RnfpAsX8hHymQ1xZDNCstqf1uzpPo5ivjW9BUzBR1HA2oBtC9
gEyJxklaE1qznW9o5Ta5A7DkePpvAFwaBybWhyPN9eodEzpvaK8RZKB2clsKKrJXZlTavuc4iWhT
qXFGCvSu7HPXyB3n5VFIDoj10KV5Ehwq6mMJ4w2Aodo1IS2RVGpWP+sJqkg0y2IepIAvgxhTdWmZ
wQdjL3IMXdatDJAKOvOF85F+bKIwFA0bwXJ+g2KU8QGXNcGbXcwuflivABbFOoDP9c+wH3FfUhmN
4MNQxAZOt/B9GU0nrXuiKbrcqsowNG6TJveOL8eLCRPqqETjoew3AFA+3j3ikx+06I/htCaJs6e5
dFSPLRJVh+UVN6ZGcZVTJZPSmTV7U08ON7sRNDpILmtD/+7C1XNDdzJvEL64cLKdMD6eq/bi3X3w
B6C634CmUWoCL+8Ab/SCiZ2O1JAFC5VsvUj559AnU8B0eXXC8fGNZKCvVdaEJ03y1yGDcE/zs3FU
Wq96RX5eDcTJAs9Fl16rK6J4WyOPqny7GEhBxANWXwJe9Y8UVYZbqEu6D972HbvaW1sqfATRE8JB
k2f4x6LCHxQhLOke4gjJ5+ZfKjxM5PipGczzyXmQFt6gl0oT5sG43NihHqz0Yn9vSAH1C10yXFsQ
3cD29c1sRozI60aCP2Gq0BgNlV6dcbY7KL9bPCesa+fsFeK5Im0IsU+yiI+XH+30Jo0Jv9hsXkSy
uhOILCd0AMoY/i68SXQNmvFAcqCiu+7Si8xJFTKgcbFyLDdtRtjiHmWh0fp1teGjaoASSGyRuy02
diV/LrbXr1RUlAE7IGfbdfck96aLLKg8o50u3TBsExXi5WsOHqYj6QFJR9yPQwr0Zbw3HPbbqqKM
fwkKJA7AgNwA4lksZZjzdA+3ttoLNENdhWW5Q8oGlWsbuUkBoYfZ0ctGCA9InJF2Dmr7VebGLe8G
d9L11RxTqvpqZ6yUkGE/3VwY1kGKu2iyjdfavVpjEBPmdrHLNhkl4bHb7Pmb0l8weRKARdIcp0OI
cd/z1Vi9fufyCieVipX0VwWP288WcyefW2lSBxY36n8EJ7tDQorb+09AEweRxmL55/sgRrQ/KKIF
C1vGl7Ijig67l4P1a6L1R/lUYlaX0c02nqTxi6ngetBl7y22e+TNXDTUdA7QcS4VFujyUtx6vgZG
jC1WaiFNRmwDOjZ8ieoXFlkjMMcXxVVfyIAWbgHZpAuF1zSd93XJJonDUmfc/hzPAU7jedTQGOYm
59v56FkTZEa0YV3GnitwpXtjo7Qp8lQJRpghkz/OGwnsDWlr+oQz+Dq94wsg0Kjpzl95CRR9yzJg
lPKxrk06ghW1Z7Qcif2j+OYSn1ZdBf704/1b9raTGwCortD2MzD36PqXvyKGYeHqiIvsm5dd6R1/
o5LiNLa5SBFvJfTV10ROMoxFY3sgeWwyMWV5QevzaP9S5SwkMQQAHeafTtDHv1Pw0+6ie8Cf2YgY
hJumn4KujIZsmg6GsocKk/p0L6hpcUyUopO5pC9fv3y6YvHoYcW5d5hN1R+0jB92APQ0DjlKgXfV
8n/3/seVxaZ/HiDPtLHLw6sVANvQu3zgua5Eimeyw7hoJDYxMpRaVVTr/eQaq5IX02cVThzBDBFz
CnDJ/7SRSm0ripddSqkc86NESk/d6HK0D/zeap2XpZm9+7P4h38BgMAVp71loSEPDanwYaC5wxNB
Bn1Zw8Bw/bpsxr/ruRPyaOUlmBWZrATj+lgdLlXoyM+nvvOZptPBIX/iEIjfyRfedVO+tmMMJTUv
5avclyIhA1aAVUz+wXbi/tzXexdCfUl1Dg9aQD4deX64bCUWBOvgBneangzhPxwzDX7lyWCvEJSA
JmqpWp6Mzsgnt1knzxabTA+j7lZvTVYp93BPVVckFcE/3+vjzv5h0gCqWyHgRtZTeMgry6L355Fd
d1SEfqxdwPVWk2pf33/ankGO1zQ8v67fxjMG+ihgzEaejWBZSgQYmay6uuD44+TzSfmy/hsaTmY7
BXyRZC4k6UsEie0O/1UytmV70TuiE6c4NBysWjmWCxQc6jCR7L7bgg8frLJr5ruH2vodzjEgD27u
nOlYrrw+TXln/UAd/3/17sCBlwnQrtGvrndzQ1VaHV5O2VVBxQwnemQQ4b2ozw4Cj8paII8OqKei
Qs2e4+JjpP1q9qEB75W4KcyxWhHTwGxm8mzQX5N5uDezJ160U4jssj89M1WF8J0oDfdWWMEUCRMa
AXfygU//kTjED1FS/BXBqwxfOyurEfi3EZhrn1a6TAbksGZZun38DqABhiyYynZvXYVaU1YUOCvk
H/cIHZAWHdoa6GZZww76RXCd1ioUKKPpTiQObvT9FMwGGt3jU0uWtT4vwMIpWsovz+DO/kOSJJUb
M5KnqNRV/yCZDjYdWJHE8qkr7ohPp/Thus8M5GXpTwxaedhyQF14WRWFNX2B4lAb8JMPm48OBfvz
+9TJ2wa0rH76kkqhZkCBJDdKekpcxfSmS5BcHwqJh6sS3YdO0ABIctUZqPGsXpivMoFnZ3w9Y1QM
zt2EdJDfd4Fvbs5cxGB1ddgrTApUsL/BK7jGe6o+SI2Iy9pu7auAYNubFrihRBzpDiozYWdijzVv
LQec9zqqcH74mpLki5EXXWASUIZKF/667oZmL94K0HnaBtJxOn4Z20UTYqwlUWQgFiOj8wA5yWhE
QLNjNBbkbYp1mhq61qG5TeKcqoBViB/bO6dBsSQ3Yx/eGpmiODXH5q5kitvbqXkg0KwAnS7eI4bT
qrmeQTn0FRi9/3kHxJos0fc79y6ZpjKaQAEELTkO8VMNlsj/JUL1rUVQ49v0vZArx1lLLurvU41Q
sXO2X8yb9G+StA/HD8P1D4SjsId21G8pgkC0t51GK4DMf2TaL/QiKjbM53tDyyzczPq5pIagUokc
wbHiZ3wU5HBzFSUsbXzL8jS4EGslts/Yovpx3LWhND1tUtp9QM67yq0Qa9n7rCcflyIkj0HPvTs4
Bc/6R+T+0j8qVrqhtV74tAAR9VbqmkD6/gLo2cYqjHO+hVDjVjfwYVLrXTRwMfFBKqVYlTOC4H5R
nqwZuW9gvVHtk4WxnpVZrY8zXJGMmO3CTqpe6Ejti9LDnnO0ImfIzhR21QMzha6zFkSQv4ZBDawG
HGoYl+AA6ePP+vpi/oO7VFIJyC1560tbgrFRLdCvyM1FoSrYdbVfNSBnaIAZrmfEN98rHw7JbVSP
lPvryeodCF61ribSMEdOHkb55X3yUytsptehqqaOEOkDnKmTcWlDJ+wOJs1PXaZcIITibuxlLMu8
X+ImJNvRpHZnAbOeQa+QoY1B/CCPkul9P70q1ueW47KruzGbVYmgYj5/RcL5ioGgEeO4GvQW1JA1
ZA2YvtDPNx3fALhHP7AmM/X35hysQWvoe9L38DP0UFxOKY+0zz4fVQicpRADl9arWhVeKK4CF05m
/HJd7CtXdu8NkFKz6cHnaGdwqN2M3snn7UYd16W/tVSGXYt5sHahOJTNSQOG0NYZo8D/ZJcOXhLN
GFSN4c5G1X4twRRknmVRGdTSZBbhrTOdAHa424lZmZGmh3XDHVCrxLfv64bmM1q/F1sWEDyEUz5l
hhBRRNY/MyLa/elinGEK8YXFt1wJkqTMSoN/VjeomKn1FNDzURw6WOQg4RDiEfWJqq/MKApkMJsh
af3wNvqWtxTtHmEdLvPYNNLPBEn1SJOZoWnHTNszrBOwO7FQ84hroE5Y4pNhp3Evr721V2a9ib3w
uQc4b8oh5H/Cjs0FLkpEURtkVsEYQ72ODaHSs+ZvX6XvL1+Y7uqklkXl0xkTHc0T6o3vb3uDm+F/
AFLsXSdYKmtbjPxxdb6U5UjDLWPT1JtPHdA9v6CD3idNshWdWzsceENVxDj5UhK5sV5dwhUeAZIY
WquBQ5alIQfeiRwkUdEyAYiQKrTHUkfYAdgTww3h0ET8PKdcC4bUFBbX2Rhe9dfTdFS+NHxM5QjT
qkDGIQe8VJ4IBY7DT1wusU6qOHZLPr7XjigRnIbnLUvbEPXLuWcwjPIbytSLhV8V6NCl2WsAWV2A
rDexbu43Qd8piDVQQrkr2JGsX+KLMw2trgqCpgl9UJU5R3AMz4RcL8t8+MQHKDru3Q0lJEKoOUf5
38ZXA/HV5u6R/wlBUnca8vTDueLsCizsntjFlHB2KGDCKZWHUcgircj/jm0aTLgV/MfKrDJdUtyC
8oPpeVvO0JIpkUyiqyLG/5gUD1uxQXflw80HBJZhK7PhOWYJXFertmuCecQwWIjuzML1SPGWOpHt
1WYwmc/u3BLVVNNH6Wjg3XeNoKwtW42pbf405B90uMX6Wwa6BN82GcBTMNjQ7E5XGAksTN3Ch4g0
A2J60XVvjNAT3Bw9Q+vWDkl+Dg1NVMnveclGK4mFRrLsovgEIygjS61Ou2tcgp+MeJcIL3aRCXIc
e+QQdUKqXA2yhP8tVlGeMnb3/RAGPLQilSYG+xslg/6DDprP7fsh1pIawT06f7RJat+s7Dg5sdCi
SsYFGZBw/67/LfrOBJMux4j2zHTd/Hqre6SyPRsimtqww9bZRmHJdAd051K6fAiHJUNjwnUKSAK8
QFKSigE+yJ1TKUrefVnYoKLjfwLnLKiwg6H+MYStUjMDxpFoo9VO9WqATcwwMfiAQ8SGSqD8o9SB
9rLYOxVTanAgHkxsq9jGJbRJP36thu8jLbpXnJYh79Si4slWTT3BvxWlLQhzAsZWB31B7vXGb6tM
8eiXxM5fkeI0M2awqT06kvZD09XzoOIjvwJChU28MpgXfSbQe6Vo/QYcqBexkTyHkzpf2IEKfezE
Gb4J9Z5wbKqmgF1VcOVMazlX0x889BMr+sMMzxIg1kYQQdl2ng0gyssD3dEeKTGeQVMPqNS0HWuZ
8uQZ3URjHOij6AKjTwlna2bziU3obI3GDOTT2rY7MGC6NP5BEj6ysIb0xnw0+JpM3JL5Jvdp82E/
/06w18gCjiOYTCh6fCbzmEvcRFM4S08MyuBF3YYfraDcWoQYVmhnbxy/u248H2nxxrDQ9YC39yZv
Zm36tjMVwptyXQiUMwUDyorqMnMqQ36tFbHwE7yEUf7qSvMdCn/xrJ940zNwkB5nb+tc8Kz9nmtP
d0fznSd5DLH1UioNwsWmFH4h7qr3Id9MWXTwBW0sPdaxxoRvZG6oNypuwDgNldgKJ3xW+0zENyLn
Oy6axuBjkEPmnCajdDJRSnw0UQn0UFx41mx99d4ThFCC/id6CThbQkhVleZp1HNhEWCcpeFhMwWP
sVPdZ8FM6f13qqY5ENW4BGTO24iuP9shVwQiN4PTPgmBOVAUETfjbo/sqSN0JT78CB2cmzBhl4vY
k9i2tAgKjEQQ62FJOI5upjYSghzO579OmKCbTOYEq9elX7gs8ha2nPiHQPZWDqY4Y6hkhXPK6ujk
ayvKRgZWCTkS3hlsQYEu7gSaSdS8mPhsXmEBji6g8/OoKsN7vD9fkMKB6a2UTrYewPktwjrxA88/
iDLaeiemB69V6Aa3Bg04IF10coSoMGEiQNQo4hYm/efr+8dkzKC3/6WsIMQygnBmFOjMzVoKFrf1
oU4rmsos/WswKxd8czuRxOy+DDdYpKrp5wHYXLa/vxeWzh2gAVr9Y9KkEn6SPkfFXqZgcIJlh6m+
YRSs8mAAJbTuT3s4iWMhnGfqYqTvFBFPzivHzl87ym/ySILA/9za83opH8v7HdrY0IpBqQpzvdjy
27LhsCcp1dgg8m48bPzO5FiwvIMrmHBwwTsY758kEW2foVrJrFJnyTl1ZhP+s4jychfyvD/AOwuz
+t8UciO88YNogxlgc+QiogtqJvl1V9Bw4GnAA+qCaSQi90EJFzX08i0yGqQxMAvvo4UM8FKX9QIL
Y10EHl8hTNwIJmE194TXzVK39sdpFzLvd551BFKktfRs6w1LnOvVod8vBlconqT9UlTZ1RxqGzcm
7UqFvJm50OOKhyzWxpSNerubEpGIDplXkKNj9r3Rqm15ovn9GWK+SgESC2+zrSmTVRuukOZLrrnm
yaldPEpo+B7HUIjdvjXQkpa0JPDaxWWMQxHIyP5pP3A0qi1fGqv7m7WBF2ID7gsYx9zzLXqeWoUn
+XY19H0U3VcUED23+gT4YQKS3zlNDitsBXJC8MaPcUAMjzQnJqIImDeAOUP5N0k1RQWfDt3IQM0F
F0o8oF8jhyRNg8J5ug04xIb3NZ9hNZP5gz963P1t6dLa6pnKAowZDeV4iVebWGSfsrKVKZxrxq0I
EqYWOJ014IrCQru4psi+OZ21uky6JnfRrnvHWe+kk21QpXD1kPR2E+HDntBTzwUZi0ob0YkvQhTC
C/jDrC243fL2rl6j5Y+4Q4m2QQZy3JVuvzZsqgfg8X5Xgw0z+CV7J87qdDI8hQ281rwu8kE0FFMG
oaM6kK+Ttkjm4375pNXf6uCJ/i0snOA9Ozm1yz4/s1SnEHNznTSFtfHqqkbIa6PldB+LIbDg4SzY
LG53Ig+MEL4pD4Rg7fCFSo65D/CB94KvaAgnY0lzLGjwfTv5bZE+ha2HA0/HHb8TF0+sMRKoWZdo
PLkNBTmHmEoWJ6Zb5R65HSMbVZjLNlAzHYhQuiDIZpp0cVVMMZwLVlBIAlZX+fPCroo0Bu3NA+G6
CLY9aisyBzmtetbpMtpj5PweINvE9RkDEWIZZKE4yy4XKJb5Xp29et7BUkhqM7tt7TFR/706jCMB
9NHkKnoyUgqj7ztQnShOjiUv+cSTXOCxDtbLsWXT+jUbAgAYE7p3hCyE+xCxrW8DVfOaANCSm26W
AKo073HoXnHZLLKt1R5eD9Dk0Wm6Xg9LcG41Sp+ZTkgc7IHwieSZcqmcy+cGwQD254MpxwBbdf4r
wq1eE0nKF8y57yDzdwUYiyfx0iqKKIp0ULKtLE91oJ4f2In+srFY70a/pAvvzakuWJCwW+5loSJ/
Ssu7S6VpvjtYajcTECcvtJkqlLaBLxjM4+T1UNCN21fdtbNSHTNqcxuXblCWfYELsiWI20KctlII
KOmF0PMlo0wDPsBLkzGSK2z3Jfl/FRXEY9IiNYRPOh/t+oA3Sb2dmfIYMHQcYFQUnWAuZnsunM8d
sYg5bYh0DrJzJjDgZJuMOxLcE/OOcKrcQWVR0O/NloGBmuIWOqZLuMF3tYjlw3rLBNk5PUlVRCml
OFLI40tEbrPgWc97hc4T0fIbKt840+fzGqgtcrpSPr+1EOENBJox3w93un2pT5dCWNFe3UZPKQqC
ob7S6BIruBEMsnKckEXGEnRcy/7l/ZhRjwosKQFE8rr8UWRAb+Fj0lJP1NPYLyM63mdItK0dbwRa
Ee23HKpOo5j9kyO5ZqSZghXTl+QZtdDfTj9JIIrSA2nlg25V3LTaF3QVXrskLBT54ax7jzBlG4gS
TrtVExaTmyCIz6pzBKYTA6hGWFbLdvCpmJhvMxrCxOT+wWbd7gK+2DF54uKjh/FmxI8FnBMcboAM
h6NcNl202S+kr7DPkblI7sWkaeIusSVBvacs7MXSUx5c4DPWGunTbQ8Ewi5wG3N6S48yNnZUi9e2
zve2l7oUKYfT8I+jJ6jZkB79/dH/+HdWuK0Teyvxt9C3Hv4yTOWlLDPq3+V5MI/aJAsmMEiNMdZ3
CluUE9spu5VOcRqP7RB9OG5KjPZtXeWQa5RwqL9eeI8uXc4OkySoRNL5Ozh1HBmnEPWCjBatGWw0
A0EpMUKQ9v++MCWTGoQHxpPk11OphvavqOp9f4a25xLkpObwbY8R5VsV4b35p43ReRp1UHy8izWR
ymBoLpWZnPPahbdfPKkYnMaZaCbtu1NXF+7vJeu0yxKhrhnCP37XmJF5MApf8rZedIlEMZOU96lG
A+tk0Uy/EQdaKfS3FWhoD7cRBoOEv418+einuVltad9JK9X4J0Y2wO2LuPqpLJ+NUMX0+WejIkef
8QarHUrKal8bfPq+WzfD9UBPBhIW7ryz0dA0Vumz8ZAFIKl99bZPQQAh9RfiqXkCYzPDb5ONOYHo
s3lfGMksUGrMT8atteQ97llhgjwlOPRreHdSSUJM7q8J1EueEEud0EuUOE8gCJK2UlzWbEFzrYGL
w4YzIll08PPJthw9pUONK33SBsVe2uEGeH8JoxTmwDYQx7xh0tcoKIEoYbIt+crUK3Z/ADOhtO98
mBOHC1DHRbIhqKySosImz7tclFDnbKknmT0f7IqXaYbk4AuBsSoGDeSVNbJFpLrq3USNiM+t/ivD
bDOd977MGAtpUi1CZ6CIy8WCNnKhsVkK8+MPvkGA9CCgZDYyzexa+QZL2b9RFOVmlqBNRBWSDI1T
AP4mznNQec+A2JtS1lGpiE2e6dWNY73Gyg6FvtwMkCMjlGF4HPjx2piWLpHI0QeYI3OF+3DW7ArU
ACNTFlETH0H3WlP3zJwEhrxPfaIcwH0Pn+7/bE2v4+YvLzV0kN5t+kEzUYm/ynGmepA83fHuC41i
OifmXkHSthOY6xSU6ejF7Y3GlME3Hrh0WKwklq4I0BmLcNIV3KBmdwiRL+xmMj6E4EFY+xomD2Tt
/WmqWOA7qf910o6YAHzefbGQ6X0IJagtPJAh3M1Tc1yfChurOnBS1VF2/LejgODbXdK5XJuqqRhd
7py70f2s6GzRl4as5ChLkkOGWcdMeS0viV7Ih9Tkj4QoCYkqPHZiUnctMwuM1OROQMogJnJ92wHT
gOF3/hQtE1N+4nGzIXx/MxoviJhQdDW6kj8NRJyR1CADPTSaFJd6UmHKv+pyjYawJjpVs//xq430
Zez0tls12+jFAcTH0ByVVblHztf14za6xWMi0uNMSZO6h5YAep5ipViYiBJ3moHw9TcQU9ba8U3E
hMl23t+b4CdPHZMFgx7MnnGv+zun2byrXOqZXItR3TXgfreaXSekehHmbEmGejwCuIS3EAPeIY9+
6kUofAsdTNb2qcoYtvazRYCtfK5CCyJyCaDtGsXr/Umx/zut+Fz3x6wz8g+75WAEUibBdHUCNDMt
1Dl9NcHy2Hjs/KVNTfNvnqZbi6KlTrLc9JLm9Y+dZEKR8NXUvl/io/ihVcqL7ZaHthGB8up8VZ8F
oMNukzHaklkIcsENhx9EhhQLgweMdm1DjABZlYKUxsj5IdAbwox9dhuL3YTecDgH2yPCieC4+dT9
CaJN1ym6/gMAeTVLinH6HaVZSFyCRfZfBRFQEcDfiN6U66wdMl5hwi5H0yKVA8KStxE1NmkuZoUC
2zjvQZLSQB+pyOrvsDYSRjRGmgUy5NTp+nHiRavIShWxYEMhaRFIl5mTiFDKJPtz1WCHTXwmrugm
DyOfvkO6DVm2jpL5q1x5KNLOI2F+AiRV0H1OtIa4ibXDh8bPGe0X/mSUW6wkW3UD8Kj8c8var4UV
RAbm+MO350UKQDYQKv9ySBGAkAYjO62jrqNSaDkV+Ckp0uepgFuEo8lyawflFpLGC88uBMldDBiC
H9aOEzHFaL+1f8DxuO33RgdKqazL4Zww7nuLCLnEWljsaJ2ipv2enNqOBlOE/JE72t+4Vg1/Ibjx
kOrU84Ux19eTrPyLZ4gNEze1TipNYfNar1y9eBgUEuPsst+P2iuWPnreHyFQKp7K8RUF9dwY87nD
AoVdZ4/H9C7ilAHPCT4dgEZGnAj/bGLo9xA3lmVMn4cc0wS7+Sp4AnMe3bayyOzfEVdKs6XuP89w
vL3UXywQf+ucuGhfNTmjCA63tv/wMywrZRRNu3NTRjizTNIUWYW9EEd0a+yO2DaRZJHAjLZgp1SP
d6wEqeeNiaX4e/sZpWN7HMMtYYRewMu5IiIw7vmV/FCt9GrWEj+MPH2frsb6nORRkYV7nhsQ96nL
uJeOUK905nvjdUqETQBMOIIQOT0T+pznhEbFx543gQG4YjxSlH8ooEUTCejyUfTpiKdjvS5TvOQx
SDKeQCmGyWcmy5TYDfxc1006w2O7jRMh69b8vbwjSDNRAvLM0e07I8Ng5CRzsVjLNNi5rofATP57
oTqqXB9ZyXoPfRekckfU3gEgPSeHPiR9nRd0zmiAjL2uew8/xNTCyzsQOj/6c5kZrgc/m5KjQb4j
hD8bNspLcAXk+oo6F9doriH3tRpZd1xSz1K7hkmO923YAELfVmK0eEGwNvsdk3h5NPUo3O+kgjH1
ONu90DuGQrF9ynj4Ej3/Q/3p1yb5HlX46/GvLBVntxfwgO3nDTerm+nVixWUbB2EajPyUR1fRfLE
romgTNjenzFagWq1m2xAGxPXP0figESoJvUWBmi6lZo4VXxjRvNzfyVV3UzuMBYT/cJBm2yGgERJ
LkLDgLp7mq1U17EI5P2K++SdKyaw8KPvCyQpDVJJhoX4SZ61NLWGo3aRK9sAlFTDHnr//Uqg30Ed
t/nNGIt7vZVBzUTnCJ/Wtpvc5hRsMzHMD8i2tyCi4oI3Ususch8PhHndXkaP7TEb/5ZxTkKCzOKs
swJwHmJrWpKrdRFIs7Wl5L1k2js/bMxESlyHPOymUsTlTP0DieevMJw4E1oTNHnuuIaXdhewZbHQ
FpGT2olTEnNm6bMLgumrADzjZcvb7hVnv4kTkq1hssp7qGoA0ehBtak0wy2U1ZRfoOxdINjuRhTD
moaXgOz2+aODezZZo0GdkxK8Z2ACP8DzSJ5e+K8rNdA+C6yCr8CA2hTRMdVAA7ubBe7aG6aobswU
pgjRoM3TOx102j0PEaiRFEw9vzsmPX8rsQQSnxdBWUKsT7Ylo+ZZL0FHXqTEcWVdOzOR6aXWpztU
gygMcdR2lv+Rc8JZiCIg2UUIU24EedoWUq79fqgg9EmeX4U+oIa5REcfZ6fHCjfYbi97SCgyej8d
cvbTIoFydHRY/L4n5xByRTX6h06aEZZt480LLRUh0quVot7M/aNdLdZGSFlURHHVSSuFxnzNZ43J
VcqXIjCArsBET4B7Y3fHUXuE/+2rx80hclPxBzqagkOCHRdjMx35TE1VeymcB2Y6gTfJRKZnQo8Q
AAVhYSkPjsfOCg73VrcDGDZUzs0w4dDf2Im9P3AlrOzr+nAU+h861waa9udrZsfdf522Ns82YXs0
t0ziYD80KSEo7GVKr4YQV92YCsmcqN+1EHa76QMnW2aeX75CJMLIixmMlbQVHpU5AoeUhf6GAETH
zP85MsDfjMcS5XbbfpGbGG8DYPsKvc2f1uMgQTLRJVPvCTzPjl/CrT87g8IASAN8xkEtCaKaJd2C
7bf7QdDaRcmv3pMam8C/NFp9+OfkATczbZb9/J7kFdvgFWVtKq2DPFLGYdjDBlgdcRy2U30BjnAj
IAEIrlQvAmK7eI7oa3z0qs2fbH8gqpBAfcUp1rFZITV7qWii6gGlKOhs/k4zXVQtaui3ae+GO3P7
A53jiIsL92AiVIdE/1wXu9JLv7mbF3enwzYoCjmYUF2j3KeSiwUW04wWFdClfJwf91cYy8NuypxE
gZkbQQ5L5qAr8T198ymw2beyEGlxHgbueJncEzGXGNGOihO8xDAFmbgfEXcVO043j3LYy18ppleG
HXejC5CcPtJEU28KHZWFoCjiCbhO8XTU7Py16gDiyItMIhmQlKcD4mvwzZYDZeIUhV/d6ovAbZDJ
h9BVvL6372h17WUK9wqYjeWg4ALuVF4kzJjLpTsiDCZj89Bnw6p1FGImCWo5ONN5g+Q2v1BuQ3Ss
PLYW4yV6u1EQTXPRVJHp0PJQqMVqT4XE+zOo4p2NPWFNb8KmzfPus7kZTYiNHYxqro97Hx4xjXgG
0MlK5pN5qE/BqR3WmGipVhBkNbKHmikOOWSS1bFANg13QEelYC85Sb2salU1CjSdCm7kR8sjD3sR
9kyocNOTZ4kSQXbc2m0e2NcMbgAznaXh/ebeBCK9uz/AlfBk2+Ex/42ad9mSIecFrYnbU1IATRxO
e7QSlIjRpQR4FMo9mhmmIrzJxRkmN0TrwVIMAJQQF6HeX1ftRa+TwlDfW2iOuKRW4pR8O4osfIJx
WuJWxZSn07y2a5k9Ub0/ksizqy919xCQnzbJ7aepUWRSq6uDq1OXQ1Ny5H+IxlSs+vxXRPqi5N9n
o4VkDIvlDS4x8cJKRJjhsDjCfWBInwuAWYc4UAqJGFyaLE9/eUw0DqSRIOLNLzASoouqu84sn+21
S+wtgWu8V3DeBhnBwoCMvZ9bBdhXnvEeYfQBZ52uN042K9ho7qmokrvDqeHIlc/kvCVeSnDk1rQt
WpAMM0QvRw2oahzSecVLI0zzYy8ufzWp8rWZ0/OJTaHv0+3XTfry0qfur5+fJ8OKpQhugd1M4+N5
m98rW/LoP2wS4k8dTOX9KshhL/Zi9g8Ij7yWWtvHJOYhZlSVspNuxVfRUd8VJHVy+iB7pnzwjDHP
dEDPGdSoCJYCD9rWH4X13/jAEpXcvCbj1oYAJBNJx8z5MTCV0IFJZ8w70ZYHpI55FJIOga8XFTb3
mdomEj1vCz+3jUFE92xEWQRpidiF9oRHPrTcCmKr3VTpP+YGFVURU1F+Dcvn2zroe1Jp94KcsVqB
kYmFEapcWNUWb/viIO/iFEmfQAjMTH+4xEkaRLhCf5Qm8rMERgS8i38MZ1xRslrVvznuuHgg7SnH
mmg6eRChuAIAV8ykTMwDtx3uepbRbUDtgFQRQW5Psf6myQMPtb1dtUOCNMkcynFdC5x/A3VkYgtZ
AFi/dYZlWeSSheN+Q/f2GnLRwdZV0QdN+UXWUmd0rN37mG3DZeiYEeTlb8BxLwcVgdwlI7Ez/FnG
484uNbj5EvEpMEZyGfNllYJxVXOnHVDn5nqEpCH3Or9yPvxGRoPC3+gdKXU2S4NjnMhvLHWcB1IQ
6BYdInBoklwKJTFIWVRZ624K+kEs4JjNwKh0kBwZ7xK1KI5//lXF40p51GE5YYeZU1G+XXNvZTJn
hXRA7efM9W5F2qBpHRveDixO8Mp5dT2mKoSSeimYgcOUCiZ2txLVUQewvSaq2pyz7XV9h3ytAUL+
1+Tba9yPZ4bNP9clGwuN+iu2sm00f5tVA1CByYxt52aO7Ku1CEdVrHtqUFboQ406hewdnocKhRm4
pfmsJ/t7H/Df1lzKEd9MEajHaQSZOYjiJw4sXtfi4ZSEVHFo1DBzB8y/9wbC8XODDbvwKQ7dPQyE
bARaqa8JtwziU7wDTbdCvTJ024RjEr9wjtvUbKDHKcHupY50n8Dfq64dCVbf2X2q3X9t5Js7rOHL
00pFGwMW8a36mf34Dnx4tzuPNZWVIDY57OEswihv4rGm8Q3LVsFmovt0Mu4QKggTnYbu4KdV7vrZ
YoZ5kZFSAN9M2Lmgos+LMgAeVuK7oyHKH9SdksRMilZu5KE/t/kTEnjeEvZ7m29pYMDIYf0vUpAq
f0YjomL274BpUjaUxipMEdfuilU8eFz6M5TrVkXh1knXjepDCWcetyYWulKY7ynLbGPnLhO2jNv+
/EuE2Zgm2q1AS6F9QRy+mbWdDNP7GukaDPyZIl3a33Ds60YDaGyYWC6YjTVPrv72mpOtUaZ0wJUh
WgnJdynyYTgl6QM8AdhKfF51bGnVhvLpiKNJvy7nBBD09FGjCQDw5CDHCYKHkAhZe8rmiIFz7rtv
+MOahBoEtuB/YQ2zauXhR7bkQd0rBOchMJ3KmxfAvxPCTwLJmplzrIITh5EQeNP84uc55Gq+B/CC
K6Pvw4wY3vyjPnNZ3rdZS44i1RtkhT5th5IBEHjaWSQ8L3SOVw6IklGCihXw1LLMrj+bAWkjQwgx
frBj4JAHShxCez0gudx0xQMGzkZc4vBwYkBuwou7go/xks17mt7deGNG7UyjSJGnfq9Gl+vVVn2v
J7x+wiG4Ru/Db5wRVQdcyqxKTMNxq/m+GLA3Qpw7HsuYfxa2JfkcjyK524NBsCxDLJusPGNjY0c8
9/skBFPrOGq0ByegRpgvHx/1d5LhbrUp4cabQrlzKMEu6KEdKxjz5U8LilY1UqlLml5W8RaPQUP7
KqJh5iQzJE2jbEfGgf4EVdra4G5EJ3EfXhtUwjhii/5qpHwfbbqTazbuwhDp11vK3bMLU+926rCd
rX68HqaAF/f7QGm9aPqyPXFA4yPnGIU8wnEIqUGPqu4b3SchqXkFnNPhhHDUodKjz02mndpZMQTg
Wvxt+fQayqCcjQG37w0wPkqn6YJWWBAuDmiYtY9x+Zul+PcPNFnpEmlBc5IKHTqNikI1U8HfjnkV
mROTtBMdtgaR1AfYCd/HqHa6VW2LwpNgzO73835IZ8VGtNa6rNqm+M/lqBT/WCksjQ3lwlXkhJbn
H8xJQXhIt5c9ENaEKawXIOnuRpL7sJibimDJXxqZVmlPAwtwO1AJ+b/hp/sXZfHw6FdaYBwW9ZaK
U0+NtcjRpMU4LF8+FbHKTEtCL7CW0UQewenc3yOpCsP89BFVmEyuVJ/LrFkK/2S9ow8J83b4szKM
AxlAXX7iW/4LXmU7QgLgS4spODyVQPa6F2zE+U2zdHa01K4kvlXCuw+kQ/nxS2OUT51YLi0m/Mvt
9fW6uE30dbjxNaR0f6qXt+QfiH+YIVdxexGj2EPFwMp3q5RXKanpAxZCXZRbb5ZlRO17p0V/4yN4
cmJjNc0pNBtCOg1vwblurEEHFoaYgUu3E6JLf1VBQKgvIEaR6/N0VFdTSfc/bICBJGT+o7joTvqd
06SDqnwkpkSmlqf0GW4SZEEeanUNDNtXGCKmvHmdjMBIEmav5vG0crwfabPu/w+MIqWYkZzYNTm5
o2Npxu4vsG9HZsCsXTiR/akDadfvb1tSVSb9KVvQggCtRBpjyzE7X28IZEQnLRkyXpe1RScVqErS
cyUsgrc+8GR4iqfh60GShIXtlPMkMJbjbKSxcrtq0jq27FMsi5QcqfpHsf0ppHfAMT+f6jDffd3U
QkhOP1HNbnsZYceCcUCc3FfD2qySjb1qUKpT7Qo8EUx7oDtbjGg5WEukC7VGYENoMI1q6KcB19C4
FqahDIWbJUeujbqox9Z95BfjsdPnevQ50GUqISWeMAbbPq0A0wpuxltrDdyfBKpQIY6FGH7ke7L7
5yR6RLnh5m72tgIzrJ0B1O/9uAVjpx9tyBOkImVoCTIHSoNWLyQmegNODh5/brgf8b9tvkr37PJ7
tRQWRXV1+WbHL5DMsKeZS7kstfA3lybUPUojDeoEgnn4LKydyoC/FijDIPtWESFKBblGUHPlw82C
TrC9opShVKbr2jFIJj3GybSd8oWTAlOC+cOYAaB0Cx7UVsJMvMWXO5TeNpm3312cKKSlHRcJISdO
3GRckWbHlCWHO4tZHnMLJlaBf6cbXgZNPvxbYl8Qnf/VgI3CUZFR7vzCvsgYm4H2KRbyNkpJ3+LA
Yoic6PbhwRCBZz0wXZnx+QK+7gh2t8uCY8PqISlzuG0UPhgXWWpOulzUuaNoNEZAGmq/oZ7yLSPS
cOT3FefArTDojOA9SafSrvBYN4T2oamzI8409jLx+/8DB9oe5fe1OKS2B4lLIrLAzJNYRsFDWKcc
fiRN8FfjY2zsfOXRpc9+XlOlMZ0b7Vq1G409A5N2S9giNAKqTsVibvi2ltSdVXxk/5tkWEVR0FzG
3h3nh95lKs37apxQOaPJr/ZdvSLkF9xgnyvPxbfGct5JPixE9SFGT7RVrXeKHdc1JFahXPPIH2T/
N8oVtNp9od1q38kY+DogGiWwefSi46w6INl9bY0HHDW8yVr/uuRIQS1nIYq8sRQ2GHp1DybciO1q
NcXdxHehJ6lPH+4GfjEGBoFK8+b3fAPxkwm9g4Az19rHHDGf/8/0w6r0WvjqpDwPdzWPn8z1EX42
o8YitSQZv7AFPpzL0aBDMREVXYgnfXSFtmZ8wMSYSA1tka36XyZutWB8qxWf2slyTgLw8qi9z7wq
12TYsLLZiFh1OiwyoyBkhZFo5/UFrBcAoeOhKLEY2RJzcfQoVn+VH9accIHCrvIKrgnjYgYVI1TS
WLzVOJqrD3EGxFiU9j/aWB3Vc8WnaByp5cIeBvatd7o03R+BAeCNvHAUHW6fOqKlSrvCd+z/vv+W
KRW6kRq1ZVtwLUMbz4O9Fay9sDH/LPrN8+jrx8Y0zjLxDMRZQrLy7SCKIlMOOMbmIh2PEn4tdevA
XB2rByptOTvQqLQbrgcQcpF23cpUCO9GoiTR8idUadhLx9ntVRGaJ3kKq8eIIXFH6LVEVjJhYrid
OecUxRg5etGsQdqYEI3EvRhuDmz1Mn0F/ohz48EcQS2tv33+6RYsRYJSkq9CbkdBC19FztDOHGdR
DBDsMM14RuMSjodgRc/2crBGMMbKxDHgVp4lwR1fYKASclUquSFC7VzmJ7OmhHyzvlFIU9JX6oZe
yqESCz6Qk07wZdmOtm3ewhFKkJi/1XVh4y8fsyRwZF6f+rnK3k9IheniSlQQJzqzrsZeLxTuXl2f
vUmk47BEjKis5xVHelBCTsYsaY8TVYip/HyijeuYrMpt1gcYMGPBu2lp+iSS7/+Wwzg4JSWkw/OI
BcnB/ncBdxwoJej4Rz6vPrVcuF/tvUyvDO1uzn/uFNeVuX2zKC2lsuSXCpEi3/vRzXCK8nfv1Vj9
D59BFRZPHF6zFxUiOooqwM6PbibPSNcxBxBikF0uSP5Sv7DDDttCnj9SZ+9iP/QuLh15bAQAa6Q3
KYgMMtXFTlB3pKmD2wNx6X0bWnRTqJgs346V8bnOLj0LQua9W7A5nJVjkpI4Hvf4ijnfp5buZZF5
woL7lgRIshItqG6T9RUAV11Y4hiBPq+6LEA64x7UYplZw9kp0Ry4B7lAhkT1EoX3QV7QVP3j4sFw
nNKVoNYBE8uQDo9BF3JTsOn1ESfXki7U63r7HQCWY2x/tMkx6F2QmyQHyFfmtli6mAWqocpTGl5z
9HqfxVZPkPqBDBu83EcISOc2YRJfLK2Cc5ofTjZKSGUHwI1B0uYGRD2zTH8FzrQk2zk1TGcxGMZg
YNggHqwg5wOGR9LHhwedv4gy7jmYpBCX0cqj+la2lq1LTO/APE9p0d3mcVoeDIHVuMujMz3geOWX
32sGhyjvVp1Z5Mlp3hssu1l0jb/MfiZL30GJT0EWhqbRT81WD9Ofh9LnCgPcVNMbbuFMo68douwY
90xU+T4lJc9RWd0kw+WOo6w1faN5aZhpRqtxlnhA4RjmTVGh70WnLsqSjwlccobBGmeWCUNLJ3Wu
JGgP13BsVznuMT1cQaYdFBMy60KyFc6E1dqQtggyO4h75WtzSk55uPag4PpUd5Zasi0ap8+Et5d7
qyPS3B328CirRDukEJ6k3zD0nF/OxaaaqQ0IqIEGcXkEB2AV+xYrlRSutf+wl/GzEkN/cpdEThg0
tmEhpnSNALDfdbt7o56Gg4Vv3KpBNbVN60jR2zLnNEHMRK01SQuIxQyKVKhB5NFvA500yRHK0zoW
Wkt30udKeuQW0JqTeW0o/sYGe/orXQL6ViIsU526WmWqfOsaLA4HKDBuuU7FdtKVLCHE5vz2r8vX
TM055O/A5pzCBbnFYBUcz3JfC4DSLRwDSV5m3oELIfV6iIEI2yLraB9k/uKtNHqdBVuil6oKypmT
fgU/Dat7mU5YcdLLOTGiZcA2Ao6gCjQVSsfkYIrjwt/HSmRqtJCnVshBbvbDk7Jh9N2+D57cPZZ9
6hkG7uv6uNt+TZnrVm83oqaAASEnLqAepjGC0B7LvkziGmNmazArmzY2C0FXGE7Q5lPXwp1qhjkC
3KYvJHjBBaXaGF5/RiALqJCt6V514JH3ivUjmnBTByZPLrj0Iqq0Y59Aszgt++315qQzm5JN/pHQ
B4iwDo4UbVhjv7rvDS2jJJ++nnik+GZPGTQDaWl4iqeJZ0aXVb5yolwjfMY/zoojfIoBDpO96vHp
C0JTwKgOW2eTNHXaamoLJa1u2xniPwkYTHaxUnx2acNZinBO5I58kQH1KXG0QwU0ZLWhp0xUmft1
s8OblGci0bllbwXEggqgxYcXzMxqDiljKmK3CneWgL+A5lZrprEVfEDMR9JfYVHjEB0jI/cZWDmB
09qwMq7oymT0VzF72yinGru2w2vDjHa31MyC2I+I6xI1BnU6wLXz+u328XsQlWRFnh6JbtIlsiIP
ay20OdyU49M6q5T11QL6l+AfFiRLYFbmr31r7OpwN8b/MItZ+SS4q0VUR09MY4kFp4OThONP1Moh
nhzpMK6ibXJSiIgLi7HaVKC/n+XqW3hEPgbt0VidPPcrzHVwwqBq1Di0Yo5CVOz+sLaE5DgFe2tX
fROgNgHiR880MQYIhd7+Bk3rYYm5wLnF6mknLlYeh6OrVevW9AwuOI+TAMcHDZK/usml3FXc96bv
6xhAM3LlOUDEZ5QJ9LAi3mQ6v9sH5m2SPlLxSRkCBxaNC1E6+OQqudXLddGUg9PFbHXsXj86WTcV
n7819wbuJYakDNBYkib6a0WaVtA4ghJ3fLVLEYlgEH9mMdbsSoUSqztJIzUcy63pGToJcFYX2Ai0
k/fuAjI1iqkZmBPpHiSMypbBrO0shXUBw16kcF/gxM2YQXn7Rox+EyFrpviusNO6e0vV3lTKSAug
jynfZ3a2vrFn/DOXIjKlmkSBZIStXouCEFUe9MbKwoAy5g6CZZu4b8zUtQokP/3cUsMRGhsWneHO
oz+uyri/W+S70HDsLIv1ttX3hZ77ENCvtYOWxtsl3r7pnsCtxgsSrstWp5K19o82XZlXOabUoC5X
ya611BtON12e5Z+b7DPZQpzhBM0vNJUJxOjbcNmTmhFpcgaS2YPtL1UM8VTOeIOX9W3ZfO7Gy4kk
B4nAHnsEsE2ZSxOIGyiFjM93hZgWLRaYitc2ub4OcCotlWgEA1A5YJ4ho41bNMGy4PqAHRkenn0/
pykV1Meq1dNEun8oJGtWmGV1Dp1Kzq8/NMQ4lnjMkVevZpcRbJUFD9v8xnpXiPZAdHM+Dkou655/
m7sjHcfSxEzRRzaQjJwy/2Ea4+0DZ6F3CNkvJ8V1VKwX8EyNgEQkm01iwLP9m7QhupQRzVLYYm5o
5MCPUNrokAaqI0IQm0X+vkZkTQ810UtDpt3IHTNFcUdXEQ+hFL2cCCadqwdbsLWV7A/RObN751cO
O03ZA89DTiGyOgtyHmEcUAZUJsK1CqbfmVCVB03iOzFDU9tJ1tb4Qn4p0l8Hy0rWuVkx+/MPwXzr
N/wtxViQ6aKUHaFHO0mNv2At5Ku+nxPPiAdI71/V4uvwVGl4isy5z1mzq/9zpik5/k9Cgwme0xD4
MUrMeR2d3Nl2iz+gjn2NSQPHtKx+0k8ZTgcj+ziMwDqHQ+cQeoOjdXmMpGHHk98cNglsk5icM5nR
0jesYsqDSP6wFAmPaf5vTi2UkA2GWV4Ymzk1KETcHwI7+nG8I4ArB6FEOyquUzEt5HktuYQULEwF
lHLAA2iTt+nQjAYgNNukSgN3JhzTxgbZCvX+cgGjZTQdRUc2EufHDrYttVyzxTpQY8c6qgDb9oio
XEyo0A2w+Vb25LfOMxs0XmAdpK1uhnObLIOvwTAk8JMbncIfMY5P4pcNjjSA0scUdyuKWsz8/rsU
rfpaB2jbPz23fVqqKhw+qheK0Au48rvTXkaKeaWsC3aV9OgAPmDUXYWlP+VDy5J7VVLQQ+zUUlRM
8Uo1AkKcbPKQYgPkGetiEM0nc/FG/tz3C3mYCY4bE1cLG1Tx8D6oeHmWpfsEjTg7JoF87uhPICTn
78pUyRJJxHLTSpEvEnXRcU7Ne1EAWpiWR5YFAqLYSOvHMoKtHFA23oYcYJUH2wtIXDjjF6RMgQVt
ZoogbFAiaTnMNtu6DcO6xrNPb1LA7xBxgOrb4bQF/wbjxZZt0iSNmnL/Q2RPcqaWo7G+Ke8XZL1B
+vH8mixfmnQ+VcqL4R6pGcH3NMOS9Mof1o7yML34s8K7Ru5eUQysola/E7O8BhCSivXwQjMs+7t9
yLGw3ivZi1DCOxooa01FA+FCGF2PNZrtKSb7+eJmLNB8OF6Dfbe8k9/hAuGbmnGWZw1ZfmwAFPsb
zEmYfk/S4snaGRBw/HKPtuq0MyVVeblkk/GHt9GeMC/lABIO25cq0J/F6nB/GAMU/Oz+K2iqX959
t4Uv5jQ3kM4mICFFRXrS7r9JMEl/Jfcml180+Ig12MDKjEEhl5fBha6aFTUz432KJf96GzxAZDlE
ek0ZUFETG+vB3Rqc1e+HQMHwk6OqN3jluTv26uHzRDIZrWtoODzW95xjXtEmpJXD9BI4f93k1W4A
qntvGZ/G5tFkXG6Uzsb9gSB/HFUFwAEhqurahpKzS9CY/5M8VTRGAKlBTxZyOEV2GifexYB6Fg+5
G8a2a2+gaDOpFu++jw/YQN+qp3lAQiF4nFIflVR/gB6WzixH4sIcg2mw/REEZqbk2f1FNlB2JdrS
Ninx86tq/5IrMHwFTpGXlVFACca2HuXzb4dknVKiAO6fSptkxlceY6K3URP4IHxHxHxbG6U2BHXY
UThhuTDIHr4u7CH0dIKzSdB7UPNqSD5iA0CsMzSBBzsNVx19HamwqrqRCwauWnFTzVxzIAHisXVm
RoahimuMS6zFWmpcodvrL71VFmSUoxS8KyFzhAk6vYWrbuOe0AsIdIliO9dKFxl7bTtFOuj965ZU
j15gBqaLuLVSw2O9LlGyqVVfc8FNLjQglzxu7q87cr5Ct7FqHbssSm2wStMSTLe7gh9LWy2xgh0C
PtmIWsa/GaUUYAvtOSJ9gINFiz6V8hGinovqni1yNe/P18GCj9OPoTD7d70tMo5oBToIGdv2fOwc
uyWwKSUNlankG4llfKUlJpJm55iCxP7tvirUbgM6/Tga5ZBPGNcgfKVqPIzjKcsqtx6NNabXhPf0
tXpfrbkLtgqjnNBiAm1EPmVb95kfO7WJKKbsFz5QCpOyauuttECPlsY9dmYh24s/tG3gL4QoeXxS
JwxPqn9EySuikhrxpGWkUL9PweBCIjcTs/OIpCX3xop0QiNfF/O8EBMeafcERvF0PB13P2zRNpQS
9ert8+zoue6pvpezJwvUcFFZueH1xTvNi4NwQqaVkHi1+hiAEClQLlGHMmXExfOl4KYR9hFULeGf
EV24bkT7p4IaoDrYCJltLEMGhutKy8kp7zZBfabkMnOj+mSB5fNftphTyoS7903+9TOGpUP6GFwn
sMjc7l4e3skv6XgU3+8a1Sde9rzQZAo3Q66ARqx8hzZsyFFncaoZxhsEg7ZZxZvhMt1Ghvduk1g0
c8fwWFRCJ9zIbJrDVU/68EH4KF2tMuqclxzFeaDDKHhmazytUZ4YJyyFouAMxSJiSlHQ5C82YmhR
317K8gdOiQieu+cHDNeVZeZZXDvNuFNCzm55nB1GgjrvMiO9xA0kanmCJfz7FLH9mMvIT7zYWIoL
ZfZczEpQN7GG3PoPPW5tThKeOdlswokFo6OKpPKDj/dHWDgh2EGKR80eeUu7DdUEasC1TJ0Jri9x
DMh+/3D6/kC/e9wtty1nxH9x9daymK8cqJKoG2N3vu8WlbY7oUUQ+6EcOQlvRRVldKBH2Jdvs8VO
HGxCiH9BrH+t6tCdPxxW00AEkrIS2qTPA8SGvwq69Bcq5hl/KJ/5g9zDzU0YY/+r5s8W2JOHWsln
j3TpoNFKNiSIy52at6A1zMQwMV+FOKvJwZk88mC+Fp/rr0sUmQ5IIBjUVEt1QWcLqlKDcRSrbhrz
MDHu+iYwzVxSjiubY77KNF8+TanflgNVNpj6bRPGMfH5P86+5ckbUQYkTmxYNWlrp155KDf3OdJB
TJFPSYm4IE9hPWXigPOBHk3DmmpML1K/dDiSCb/tHH0YgHIrot+ML87H+UQ5bLxnF3qzqClS5Hxb
X1lEbj6qTFpN3tiLT0c/x3TbzmxCNbNe1kPRRpIcPQRO9Nc1do8vdx/MXlPVtmm2p635kJlPoL8q
8X/Q/bPFmObwwI2SvMvRCA4vchYb+33TeZoIwDsWVvm1tpRpZQTjue0//H+56Xx2AJI05+VfCSip
MnjmcWiBbO7x11rPDSlwOf0jizcH7Vp64qWqwGHKVB/d72owGKwS3wuJVhdl2Ic4XZp4e9d6hf1Q
tvjXGYEXIR+xc9bmBaxBWTWwsaL+rSZ49ihiFbXaJsY38Rr8cPuO1SsL8eEE6yW2fG7vP1OTHF96
/wkQQHXEvDla3vr+JWfJlbNYTncgB2hQj0MdIKu9HCEUHGk1Qdw7ztxLtDLpeRbkdn7Qem6pp2Fr
9XtuDZWf7Ao6e9gyZCjd0n94abHYMxz0IeQ+gs2Nsuyyxk5PyTNF2jw4Z0RXem0f1xrH1agyBbg8
bcC31iiixw/7mM425Fl9TxEpNyRZA/Chm70kLV0HnxwPATu+3VNFsplMZ9k99UWBeSz0KoY99Ocl
N83xcPqBAr31Eh5AOFFpQg9b1AlBs6XDbv9xYuMrbmmVgJ3BGLfJu/IobUx4Dc1AqloqwLcTkwk1
JQ4sS6LhwzQaXI+qWzgpcNqyPAop9e+sJPKGKP0OO6Wkruu3xnOS+wAM3BhOTuNAvHKv3uaIUbAl
O8Fa/pvaug7ou9E5lh6+sx2A++XdOc0yeQmmsqPXEpICTU0CMCBt1dvVNcCZ7GobAqoOI0SKKAyn
PFzMM8QdXXTaHPMPyAIYVwmQMDh+bs0TnD0PcwfOab7atAHgkSKH7h+wuBHyuiTLLR1G2yB6oJ82
6pQH2Hm6WVEsBJTa4ucjsc1CySTkETXlnmS13KiL6F+f2NvAkgvP1urnH4/xWf8Jb1uQt0NlY/YL
sHWnNzT4WOJYsp2sQnosfsZymPaJ1bmDZY5tzVrim5cTuOMVLg7QNEF8uf2lwKsl4r7XXBoNKdle
yaX1poY7iZXDMCftOiNhlkNPxhnP1hf7Fi+07vZTeUdI54/CipGlcCJo6ZfCnQoNhK4wKp8a0hIC
cei8mY6Gg5FGnS6TOzkLI2U1DMac2qfGxNjjf/e1n9XXJUxEDsxW+YAvQsVilLn1YPC6ce4uViya
G+Gu4T9TdfMEl25wcCGCCWdKluFm9BUtgehxMNeAQ/9XrPdX6BWAa0advgyI1dDoIHJgcYCkpllH
cYx7pEw9EumfpkkW6X0FyGn1YO/pMPngvojnTkzKLwHu1aZxQ2ygz3pqRXJ/0VCAqR51jvy0TubI
/7gC90L2YD1PDdh55KFDCsNE9maXAHHC5jTaDIFPecP2zJvqiwP0ZmOQLNo8KA6pjKNZXhohiGWI
zEOV+I2AIQluKbcq6C281ur8M4M8K0Z/SYJfbVkWpipL0fJoZVBRtUPE9Qpag0iFhnFJdhuXRAGp
MD1Qgj1Gk7LqBd+Tv2UYME0zuRx7QxiAVNS7o7ElhSMg3fM9h6PAbPdydq0hKT1ssOSg5JEvxTlk
v6tJeg4uMR+yPD5GokprhBr8eHTZjchz5Qehp7ZY7RpvW7Tp0e8L9DJR2M9QHfmOjCFn36oQ3i18
c75b29xFkhINajM4LCds0YH8vybFH98ArfY8js5O57Q5cMdzJRchgtfzzATIaYKKWZq/3/PPJ6Ui
BMAOI8XMxuu21FxYrrM6AxzSp+BnDqsznycmz0n5M7HHP+qnvILoo4Heu91qkpEL5bCTRIgatSWC
NuOSI0Djl65OekU8MRdX47moApl2IXTd6gpedSZfmqHU+7lVAjHdeLu4vWpO6krT2LuUgfcUoxVg
ZxjT7q8nURFcCmii/mzsEml9t9xZOP4VtpZLDTVra9MCIDPUGUVLmJHdohzE6lNrHAOPmsuEHXvV
ZdCeIX/d0Aywb8tXPoU2inpRCRlNCcFDu+qnh1Achij+F+CYVV2XHLywNJmAuSlSuPn/1m4wBRo6
jom85oPrmnNXilaAFRMbp9DsXNueeJ0b1LZEoYDsExw/5SjYsHYTzF23HqTnWThRAd8T6mNpmlfl
9qE9ojlPKWUuHGb5+qt0XxLT9xrHd2RcVE4LfReIslS9zJ3PLvd7U+ix2r6QQPDY/Itj4XpEDn3l
oEnQLX35UFlKRfgjcbRgdLukYbESSpQvDUXknBaWIPwP7XZISoOSp81OKfK2cyzo+GHEXNlGtCwm
7VgP4UMlQS9nv/7bGHBncQEpZ/jYiNZBWFlerawd0MnPOXShhT8Co9mXT94fJXFbdFa6NDDevI8q
V8WtoydkxzKr/0tx56vByuFsIZ05C5/nsOtvCkzAdwzPJEIn32v/NOB4qe7Fqw4kNQMPmWxAF38z
y+bfz4Gv2BIFOQNMtqnfWlSiUSsRHUoXakG6CfYInMaJJ/fYPtJMBHng/xUDj35HVQDRlOPEkonD
iuJCVnbLXxa/C7CNnc2EizO1vUYw7TkWl7lCYRgZKLv2rHH9tFAFskdoEIqFQMqqZnJt6FBzIt7z
SI+WLRlG9/OXvtMELZjOPNma1i/rTwWqnGm8Ot4wBpEd2nRJG7qIItWzVewrFEQ+8995hNYCiPiU
HjmYcgGkp+WL6UZ4wNcgNjPeXOkj3fFQ3+fZv6R4raGkNvU5QI18aD/BIlBLFeyo1o+wRhlR2ome
h9Htiyg6mwzXQclPcs2RSW5NPwos6gXlA15j469rmv5gmUVprT6QUFNx4sXQFG9XoJnUptmosH62
MLTuUWl1D+MAl56fH64v4b+XIQiCOzlnl7+5CFa1lTk4XUXxU5tktFEXATXTTDpfSDFZd2f0ScFm
oy/igufVpb+HWgDGIGV7R7HjsXgm5A/ZOJq4Hz6UzD05qajXZsvN3j3LZHj9CFcUVGzvTvxeB0m+
7Izep/Nz022c9Pc+8w2W5Y9Zdv5kviC1MXz0Di0IpRctWnolVR3mnRSMUiJo6HpzrLhaYiGwgTBI
vds11tQXrgS2okjwfIswbOD1i1vXS+H1jBsH2unaG7iV0zbgV66KczkWVoRBPtFe+yz58ewLgiup
V3TzoanhfRC4shauU72IdK5CdfH9dd0qcBQ1XNTPIGkoJgH++tG4Ay8zeQ+I3K+neNXS2ufk7xEJ
bVy0cqmSKEnenzPtRwpntGV4CnmYuHuyCGrQJgpB5xSjSvsWtRZesZU95LAZZwFZE7VShq6Pofnq
HLEN0vyVc16F1zyhR0YjB5/8rNw6FPMZDtkx2XUNlbLnI1OKmijflczePU0OdOy126+HJ0ULVDkj
1MpeKQRidZIiPR81Lsv9s71LfKAJEKfi8x1zIUoSpzkkPNyqUk33Eb05sBAVBpywALrd8CrAlm1O
HkzSHU6tBdrq3aRrP+4PHsOx8JAaA3/cfoWEliPRdNAmL+BWuyvFOmX8JurhrqJ+dcxPcJ/L9UNt
nNlcrdpiczlcSknLdbVvqdPN1Jm2u2wSFChGYb3039qvDUvGXgJrgdG2gBt1uIhPpJ8kb4egyuc4
P78TE8QM460p0zrFY7v08M8BuqU2GFJsrcEG1rZOo6GNa1sQiaLGzmVOHleOeenfjYGL6oOWgR9j
+DjOMqvxSbsQsxgKZPUTVg2lDw/dY5Yv9pE2nOe6hnylK1Kl1e4GZVYi2UWAtUa6uk/xLdb7mF84
JWhyHLfaKLuC5IXuPZjOuFdcoAw8Mz4wYgaoql6ICfH4yhifbjPULX3i6LmReWkUAidjM8UlP1T9
DdGsoW2JKPnWHRYJfWBh+6D0MnmlndZCRMa36P30q1DUohhyyybnlBtWtvs/DAOoqWkJeZyWJTdP
NAhBszVLQQifxax07Qptz7y1jNkwXgC2tQEaqBcBrTHv5onLgyWs6KAPB6MsRyM0V0PhPsJfs327
/kAeBQxR6YoQ/9xpGLOG69vo92D0f2HEPeRsshoJvTeyoXBWQUmtm73dcsT4/7ERon1raw4N1jmm
XTlw+RuY+k4IRc7WnfwaoBNjowrn/Jp2Q3xIG92zJSmxbnMmiGQnxCcDqATmuLmHhi9mSIVzUtPh
LpAJl6wCPA+yZjtH+9VPhtQ1r6BArF72tC2W/IADYfIDw1qP0+YhpqLNJ9HQIfkCbGEWcMmsrHfa
/VPoK0SQEWt4h3f40IKdNGsKF1UKU8Exxe/oMKfJbMLsUPvbz+fZ6OAkG9YNUAY4cOFYCOqn/uuW
hGDlVAtPbk/uPumgtX8dQUMUZyWnBGavYd8vPP6HeCCKl7Z4FScBEcsNEvcIY4gMetcMTwni0b2o
mUpC3HCiQz1wgIzubRq7N9QPF5NfMmvNui8tpVkJGG3LCCZHBUfNL/wYjQ9WRxgyCGOhWBf2iRWw
bnPWLR/wKBlSA9mt8sdIEcpCj9fkpGJqTnQ2UzPG3IIw3IcWOdQxGzVq10g1rYgfjVutehlYiDqU
0q42V8LtxJGyU9hnx/seGW3UR6TNe7EOUJBB+d191Jij6DUYJjRDponNAT74LXv6QT/G0bkeuUws
LnGZTrsIRd7Rj/IW4Obca+Z6+UjPCK35M0MkKZy5d8/yMkAjLtAnNPmH/HemhmVaes/IayWV1c8T
Ao27Uj2rPOokcOHZP2Q/3qWnVQpDdy5LcicqREHVTOY3bQM3GHhqRzX3CqoDCmeQsKpJwk8nsI+b
C72K2o7FhSId+rxu7I7hwQjmU5wWpMvDov/i3WOi5XdpNoeXBbt90GTFLLm+U79AqBvXmBOIefUy
u5ChYiI9TmaapkY+qaeWNE7rrM5OpnwhmGtVDkTOAfKRiHZ665eMetMSew3pJvQ3jYj7UUwIbeSN
EYwp7cLQpQXhKX5I+uZ5SN5Zkkx0P12HFiPHegPlFGWh9cDxl0SqNdLHy3NSKd18JC3XLgpEQDng
48lQYlZkoJRhlcYFgVzVtBO7+8Lu1IZK9EmMbsiXUOaZilAlmNaUXs0jTm6L+Y3KYK50oP1LSPrI
wYO45W92gWGJQrWBm5eEu15owXF49tp6FNcsCyJ+8ud9BsrkxNk+ZsuLzof3ydyNhBAQNq9Z4Ige
8gyL8MEgTQETvZA5m2sWZkQHtk1PAZiAL71tl+6fJC+A/yH562KPR/qSI1eaOYBp4gcuqTUPSysA
JF3s5dQJsCkgUfR2qvuIcqjgfryugSp7kglGM9pV+jkEMpnwe6R822u94NAphwuPlitQbhxChxkK
fo7KETa5HKwhoJWsO0A1PmhGdMHOsYXssiqzz2gl+S67EGl4oJnxTYarEkp2YRpLuHHTE78aHPkX
oUUiwuUefpQD8rZpPxIv7AuH++M6bC9Y3Y0FzHnx7i5Qmh3Xpo3fiMwxOctgtSHpNTOXnI9Nj0HI
orFYNTyqQQkoBrL8gPUvO1YHfxfEk9qtiW+OZxi4mhQ6QWLtBtvRlhB5EQq01WavWHqRAfjr7ZHc
aXtV1OQbQvRW7SOFPFCzkrgKDUDqTCHo9v8q3PLCWCN3BDPXxryOZOV3JpAjR44sOaIdqzUc437+
YJsg6lAiGWVIdNcYWbijsgFyh6E/+nSFs181nXZGJcibOnrVGlNg3lEesCmE4U6vU5HYuIoo8pS+
kGLYf+WLTFCDxZGf2mp2IYmIcug0BPzOFskBpVHfdwMGMsCuhH7Edyu5kt2MRhJQI22sC0WUInxC
rMbAdVZbYxBgLgUTiFuqrjFTFyFvC/bOLA6C/XQYUKm6ktVSN5aE/xRSdxb/Kc35K7cLdjRpXaAF
OiWKV0ypxQ67feBb1plB1ck82Cc2VFJOyx0f7eo42SSacVlcFhGVZTOE447O1Aiy3dDUi/13a4Ty
/2jhsJ3RYiR2vAwQen8ZF+E7ft/v0jSpi7dyva9B3JZg4sRa8dQJ4jzMeEA90/wnB0rSPDGEOnAQ
x9ffYMeHis/ASHiV5S/Uu961eATt2/47RW7GH1Lgr1lMFwJesgK28KJ0tVQ9t3l9n7EfwHt2XuOn
DcmkbzPohiuJRF/PLTmQh6tsulRPqmNfcreU5kms4j4qiaQfReEFfqbxe4eiDJ+geynske7FiQ+x
DyXKMPZ/Q5EoDRvU3PRS1en3pKQqw6TpnLC6uFzC/0iDA+GSj1RM4plewMPqKILowqJ4d0kU5KuB
0CHWKdt4eQ/8UAqjJr6E2y/8pV0kvfurGDTSzaaX6CGSQrdB4j+BMNKmAniP9Rye0T+bqddUmSJR
Y7x6g6zVcHVti7QM+pAAFfCprh6OzvonAaw5pAKCsyLCJCvenQxGRhkP4R+hBWhO7ohvQmZV6DUa
RLlMMWXsbUki4uzfEOPTSCoab2nk8P1hQPBT/dDhSkLivm3mI79TGvmvCPSu9t8+XC5yTkKbi3hr
EUJmoy6aCUeGO/KH7AKxIqOb9336xWia+W0pdCdwztxXi4XA1l+MIdOtTz//z9btQYD454mKyZoG
t9P+bbZL1lYRS0//97obgLj8hc3dGDoYBP7pGRSzgKtbzcnOdTO3vhLtPI4fTxE/hKqkZd5D6uIm
G47NtfS4CZ1KxiN22m/BH7kJHCUd9N4cKnClM92/lFsaYPFY70NwtldiM6d0Y+0D9XHXH7gcm5H3
JeAOZOAkD+vePDUd4lbIMdayA1FdFObp7BrjYNdJPybOryMaJK/pQpV2eqTba0WWf1Qbcg2uSP99
0mrejX+iUqFS9HF70GZ1fi10A8ZQZxmroGg93f1FTXFnCRAJO/Aom5YFNg7AhEVFgs5c7dFSnEQn
RuV7Zp2QF5KkviaNrIKw9xoxsawOFbSoo/P/lF4PZfTqyQxJdfueZByisXKhxrtQ+AgkZkv4bKhl
zUZEmE8AUnzZLoMPPqxRJalf6p21Dus7vXTkekx9vUUKNq3Rm28eoxad0Sx+Go82FNuu9ybWozfi
cbpFcCfHNtYHnReY1pNsfSbpGcc2NykKkG8iUmDZnZYPMcVjTb1YtLHQ/BLu60YPJXHNQ+IuOwi0
NjkwyRIw8JTb0sMXZwMrlgCbMZMTqGX2/UIBBdsi6YOkef9ZvHvBgQ9cXcLrhjvSVinR8SExAaz8
/Dbx+3Hx0TFQL71ENyg3yJPC3EfCU/KI1PgwOkRqfOQi0h41T0j7DdEx4ty52osJf6SbnfuelmLu
cd4bTlq+WPDnDkNQfEwz+5DQ7i1+Hprn99lPT1XUzzeIIFttyw6njTdreAeAyxl6wLLV5vV8aeeE
tCcSC6B7vi+Nfk0yu+uoeHTwkLEtqLGrLne6SWqVt2H/q24SnVRWL5ymoQ99kKUXO3EzxYdSb6vf
3+qDYSrp+c34tWWhp9g6VPGDsI7Ny462REQ6GueVUJ233AdNbYVmiUKuM7pYfUTynSFC3jaOdt7w
M1ZpCvKsEPGGhkcU9tW0r6ATJ+9dyCrjMHQBLxQVnW4NjBryDKD7215vdnvpxP0elqCKX5Z4iEZW
xVc31JLAMxBOIzuWQm6ecO6FvKr4RrzmIzRTyW7yUPF0xgFyBsjWLEw+U89ZMgJQxv+MuHSS1xxX
zlPjF7g87ZVVzbBjtPUHSajMywRTAoM5QwebriDfWGGyr9L8TZiOrkG0eb0EJWwOuLvf3jsJEeTK
HmlBTSIOT9QxqCskjWGhyAO/6NKH5iEwZXiEtTIj3TPnca1+j8ATPZGz9oEpPQjjWDFfMChVfFEm
/wjBnA7uPhu4UpwAm3o+Sb0jrkaDtToNaTAbEAH79bCDLifX6eaEINyM7j+aspHSpjCbOaNW4bL3
M1Yoh3q5Q76sd9LSj8mdMo1cs/9Z2zybJmsL7EGCnQcXOnlkoDTLlDGflXVdA3mV1UIYtLsyqUYz
yKeoeoX0IX0tJAzznqBG8s+LnJ38CLkTKTxPxoJMgMqS7NfQqabl8pIs3uX8FMmJR969sB+Kunpr
sf5+eZSPNsfI6kAiBk8o8mYoNyo/N4oqH7fE95MkJ7rzKvm7u8dIALsTJIt1pC+Xdo7E08DaIoUO
NXRlXP59IQ3F0Y27d8qo9GqrdrarEnlHSwS8PaFwhNIxFaDfP2SZ25Z0IsIhKO6vvXFUjm+mLNgI
1eLi6IFjLpJU7MRO1nKERs8LQG7V/6Y0P0O6GygvMOWzennHIIWvoSuEYMtXaigSY+SezfdSM++3
+mDCeGucWWN/OdUEgDrm+E3bjyflzyysx4LgQQQkDaeb34In9XvLqc6k+mZjVW9px2gFsBSZtzoe
6zOfK2FwTZuD8ohQ3MGesPh+0YvtwlR/9hH9XyxHN6Fxvk7Dq1ZTzcmufXH6DRu92jdSFcOjL0cd
GYvQu2TU3+uLXeOlxHDYcXksuy8X0Rr/vPEORGMtjiP16GdPCVDGzmeDvOTwIJztOYHQMf4i7vo/
hbm6w+G0dNqRT0cODB2o6nY2MDJRkogpEbEBHyTU15w4J7HWR385nzrJks6NMJVM77h8Y8xbySUW
DZdkf+5zTfQjCHnGFS7CrJJQyhM+7V0Oj/asQPMY+CpVRQbv2OHqekGwHC/PZpc2ST9Ifcp6B4BA
3vtn7McMUJa/CUJ8wtMhNYLjN+ZYBhnX9zwlb7F+UrDY7KiMjcY5VjPMkBFTuiwUXo14/a2k0wyZ
CkPSDvCRg6u6fJqHosGPLWqaL2Lvlp0Knl3uodcVB7iUXfgeCjrtJmcnpOD4d1uXCZd8sMz1Mqqf
QGOwXWDAUocXx3ZDQsyaZRp4y3i64rDWq1Wr2qEnZsK8pBJezAWjwHANz7ZRcOxwxH3nu8di4wlE
sXfB63VlI6Jq1qwqyG740JPBUQlszgqU/QOYO06d11XdOUAmRYucZRryOOS6qS5BUUaMK79rKpWQ
kl6edjyb0bx1YtOQHRugxa0FiSJT5p76Xv+Ca4RFjxl9k56mpFkd8f3tzUK4sZHJqzshknzFbUc1
91aPZ6cMjD2e6TJw31chBT0Zx2agkDhRZNIMmE+XXGP4Q2cdbtzirJzPawDxj0Eah+665Yy5/adL
lI26Aix+MgM1KHM/UFUpKjj6cPwjEkGpBHyWENd4/XSCDYaSENgpsUxJMDkwVyENRIrU3bL/JQs6
9hPBK4Xp+dZMhG5MFKGj+T8/LYqaDFOsU2iqLrrsQvDWJjZrSWzKwE/M+15voCccGPWWVRIXi8e8
BbXsAUzxomLbaVBiQxwBPsk5Zatl+VNnjgmWAmJyuMDuqyWcAlIyiptWAQcAOhZSAhTvlD92wVKO
Z52wZ7Rr98qi7kGZOE3Y7PL4h+yAR4g1Dks3nmM+odZ03GWQchbhioza3jwtC+u1TK5w/OWrAI9S
vXMTr29vbRXJiX4TDZYyHTmHHXEo2kXDWxCFinLRjnQcneVtmY/O7iPooDHWjWAt3cadrCvh9pMJ
lUG37qpDUHNkT4FAhC4h9Bwi/KQF0nyl0eJ09Y1rVPZ97PquQL38ZY2u3HC11gW5qWvOipwin9PK
K5bBeQ0g+dGjnyMU8x4pL6rg+zPu7213ImKGEN1XGzUnBgS18Q6c5q4vZQETh4SfEUv2Xi00t7kY
fZLaFjC3zkFzUXhOmaumQz6WT46/uwzeMJooRgKDL2iqXIYt+sVVJLNh/COkGwaZc3N83cq22p4O
7xs/TSC5y7ybSYW/QBg6P2gvAULDAA8OFwZjlalAy5kVD3FfDm5dr3t6yTaYFlV/hmbLt88POqFK
R3AxDSdracyi8C0HX+vgQz80M6anTHbtiSgNagdDO8fMf1ykYUxywZkD2nVK9RNoUkkRGDW9jivX
DTuCrusGcEr9S46bNluJhbMtrnfM8Tb5CswFIbaf5T3Tsu3hep1PL/1VQcRpWV+crYODPcZbXuT3
91fnzGGKRyMPuv+0nuF2Xof8HBRRSHNuMPHpNCyUSB3p7D2w+LgB3vh9eeAC0mUhhSJeuXZgg5Ez
r65T2YFxeCMWtpZDyKoKflBZa97vPkH12Ahe4lMCeHhfgvuy1UBLpfWopu9cgKtRvvLcuDTVuz+l
A+3HwoJ0YPjRKTHCuSFrp2lEeEzYeIJuJAT5OWg4fIXlzdR/hxiOH85BAVzPm+kPCAfv5EiAumz1
qNvPDgnJFQYcLGLnnYnk3y5YTilTmVHcI1pFjlV7vuDPvOnG15Evs2qIRrYDS3B5RXjXHc1grVKE
jLSgNvdrX3qy3u99rVwcYHkE9+iiCvMmf3lisJyiVM5jzPLkMz+T/yzXE4Uj7HP8GhWZgiP2EIw3
q83Bht9wORDApP859QT+CJFdLreCjp4mga/lszUpDtIUc0xS4Vz93TFqrJomNOn4bLfV4AEYmnte
jD9wn7XBqxt5inz8pYcWfxa73b37SNptP7/h+btixbnJpJCSxFQdvdV34i4mcwa3OkRcFwvArcVk
uc4juW+nS3A2OlcrhxNJSL3wOa1f5QGNJ2WSH8HP3vV0zmACyuvgT1U5VDa+x9SpjPkGUaUBbDNw
Fra7k4YygcObMvjOZKcdlHRnOmUfUYOMJ4KTqStEFm+XphJ72Scwx9iTZe6vzn+STlDrJqemT991
G+jQcFqwv69Z+Re/48JNJAVpXWrKJ8PYlX44lGjPVoI1kp3hb0hhh/DxFQeYCCTs3UkG6XdmBJat
EEwqDUVbubqR6dPF0K2pqkpt7avjL7NMUFMBlQErNPzdqfFEbiM3JGzYq5Dz63AAcczxlV12ggPZ
eoY/ISJzbmzNq1LQNFcNwCt2xTqHFuu8qmhuI2T6pISSSbFkaPtVki1XEZ1KR+x2qDEuwPcALIo2
V4ZoNuurNXbUx4K+1C+RV39tg6zddoM7xSy+5JarrK5u0ZuGKhcZJ1LI9yRSbVkyDNc+zETkvteT
qustJ83L6JOI27VrMEvSJhcE6ira215tdoj1Rd363Kes+LELqP9phOZDweOWoVgnAxTqd+789mN5
sfYTBiILVre0ul/VkTVANaVKBjWX+rYfIm2HId96u5fqcn9VxlClVVMBfBv25foNDBAshc9DkQmK
d64/PFhQ32DoC0bqFSsEasxaGNIUUwAMyJcJpD0ZKkIKVi5qBmGUpTIB4MJxMs5lQEPHn443nQw1
JtKnO5gr1T+/MNH1LMsLwq7XAZIH8V6DYB/UIa6oiUF8Q3OoESJ7hf843rh7JRQ9BDGiLMJHA8mp
L/BZ4kWRsFpzEK4TSF84vxwgdr7x+GASTdWhlx849IviOXTe5vtaUxNiil5y03L/jIRuWZR1xqyu
uE2PU3iG4iIXfme3U8Hu4b6wq9CTy5swY1uJ+UCQfj7ocJslvMPFQPz+Qr/Fio9hhS8bcfzplFZv
wa67JSVvqJPGzVxFoJrlPZAoJw5XRQvBSptCaBUuZHhuzvEYahkbH+gaFAhbkb1Jvs4qqmKbUiyf
eUuG4HaTO9A71wD1jWZTihku/Oq6ha72gNjFpffNLgrFqWfC4ofk1kufyi4GoR0UKdOjxyPhJZ6K
4sz2ld9zZhGZsdO8se/1NSiHQinYxHjaJu6M6vThxzm3konwzi0Jk9spQIfVSuGHwikOupQLi0Kz
jjKXEqGbxt1UbVFg2ze+cY8ySh/jcuAMaGndtQ6e4njOXLp7moYll5Swy61krAXQP5SC/UXF3Rfe
ky1E7BtNhxLpjECYSOkY6gQuGubjsj+giQuFRselucNWiNcsuUFBnNxFMunjyfkZPwyA0NUFLmWg
1uJlK0zsueWu4wp8qUfwdHOK3gJtMnKQU0Qud8MsBeqqNHspETvDd46NADqPpWSwkL4KR9clnPjw
jaajuQ0Mkvh43yRiy1oDd/JXEADe0vfRDp0ei5/lq7QTY9GxrJPOf6J2mwTw3UyIgau8tz9F2B9P
wFayjBw3HAxxftQlDZZX5jiqxGhEkhbvw0Wd2Qe2Ia8fZYN5duHoi9bQ8s6aedOs+su1i0Uvx4gK
+i8jg/HmRHRfla6XZmOAmQgd87pHcB4yu/IQvvtUxotndejOrbeFHudRveOx8cDCsM+5qyMPGkMU
06MxGwPxylkmIGU2Y9ciijZzrmLJfaJECBUu/gJHd1BLvMqD/xORN5I0Kt3segwa0Uo9NcVCktGK
35zp2xS4t3a/DNCyZDrHM31l5nNrHoDUir/a5PoSxqvVQR5PtmU3BWXIcCuK41uM0qPStW1PkBwN
uTFD+uhUP1O1cDhMdBxGnO1CFxT2Cgdoq0iSvxGTPSGRTwFULb9r8nNp+NVK7dC8do2qosPGVrfx
QsVUS3ZqYRtlxV73x8RXtqPGckXAgYjb+cqJA+Ng49oinYi/pMy9SFPnp7iWexFgxhJ12VAAX+PZ
8ItzRwwsB9LaDkO/0UuwZ25XX7x7qmuMiq/mXuSgsZJjnexfH/u5s2YYB0xlesXI2S3mmd9yOuPo
znOgnSSGnFzFwcCjzI6iVIovrjib8Y1DcSjku6LNSjkWYfHeI1HTZ17gQlYq5Chsx8J7+NyY3IEc
Ey4V8NmC8hzbO8A1saLCQU9Uwpc3ur0aXnSi/xEXau0qTVU7pHh6l/rlVV4bMMhiwaEeKsGUusTs
XLcKr57myQbIpAHo4j63ss8tRSYvfgOurg7PAWUjzpTGIXGvXJuJZKqVy+I3IZFtOcAhW82fdUNr
JRsQlKRpjXfHuagVU7wBL2T6/u+KqySfsPG8JYC2/SDVNl0tdagmbaJJWwDEcuwren806fKxHTJH
qpaJ8nUQccemjtV+hlwV6HOphTplmTco+okE9VnFGLgQvrNl/OOWBT6jffVL7TcrRfLHbPylbg/d
NMnmhJyB5dKe7+NJ/3IuSiuR417CoHuZhFGBzD6/ubGoLkNn0bRGFuXFDQQ79obKnCbFzNFv9AQC
aLwMWzW+4l0ALPM/M+qpVGaFvu8s2TsG55K3lRn/cS666wH1N4b+XgkT1cC2DhqhqZKm4fPLyHOp
NqJ4DsDAgPRrAAi3Yvben91sS/Eu/S5qNagjj1zs8Tu/m7eHpG+p50Lt4oHmm+16zUKzMxJ7K0SP
QC8yqF0Jrh37YJhS4CGcLdSo6D7XbJIyDYj9VckDggwbkLn4QEnpthQIAxMZqFgd4dE0bNZXkxOO
qOCx/0iN5XO1KVs+Jar8j5CpZSOgbY75s/n873mpWjmMeHIqsYD8fT8hWSmc7B0Ca5CLay5HzplJ
ksegX1h9XEtNxeWztCapGtJ870f5Vl8cLyWytDEjnKlxQ7XWZ+EJzCl/zNBYho0UhxsmSTtzuD8k
1XLNOce0D3YheIoyApSWdAj+SlfYCLBfETA0mKfG8vrH/6LnAIjbnYYTpfHMlOTFFB79YWWTVwnl
QwjuhoW7/YqMSyWaIC3YYpn9/R/X4Wa6a1d2DvlGRxGZTSh/t6pU6TzZPei+/v6XX23qoXzPPp3x
hjuMSWe8pcGI0CT/Ldak2xOtUz6NDcdRoeheAMkX/4lfhR2QGEM+DaEqpeugh2N3IezL46isaTMB
x8JI0is71YsIbxn1FlBu7gBWGiNYT5jmhETL5JRX2e3BoHu2qC3v/4nCb41bv57qVz4SWjBXXYBs
pilb+p642PH+ElfGzOHD3ST3p5WyAaX/qxwmL0cTRs/yDyyHJSsj/EosXKrm10ufMLUQ/ATh+hJI
GVtikBOgRhMZkC1yLGcsaoIvXMojLxwCgIRfJ7c77q5jr1J/vt57E9l0c0LtnQYkiX4cS9jHaEmC
WSgCkbAcsOWqc/ey7LqTAtuXF+9OFic/Ce2EgwYkdnD2dloLmSPYlwQe0I/+csvZmEVgaUau62c2
O7loMCSjShezZvs2doL4KBxb1ijgcr3Ld3EbmYfvZG30sCvGZa4pLn5CL7/A/vOx3uRgP91jWUZ5
/QxUphZLvfwo7UQ+/lIBnEjslz3OsB+J7PcMg43NKeLYsPDT6E2HfTakh7WG2jAe5rvBK9mjrSGo
e9wIGhF4sVQmWYtdq8ozjldkfrSu99YehDYSKdK0uCfM8+h9GjYTHE1d39Nm7QZVaHHGGFPjjHhR
bsHCdgJ1r6vPJXJNH4wsLUH08GjTkOhVzBtYdMHHoWJGenXOSKbbaaSte/scypT3enWtSQRiPzNi
SXJO6zsN7wcLZs8VxKUapMNUgn4/gwWHEKHcsl5btFPQqyIgbN9urAIpQJkinHZ1Lm5qlMLbLRNf
75z7oPSCHYSlCyNKf4JqD14zJlc1723tcxdpIstqlqFdinmor9JNL2sNAUO1i8ysg7Ifnm4Vgb+n
kb8iz0voZyUHWEKQfpcYziv+DVyuDCoLEPgDSp5e6WhNmIt36jCuOEsEFdGF/tt1WChStMkDOUg0
xZFr8fM8Yp+IWt1qGtoSG9pFWsMz2Ux5qL3pmBX3+mTgfgmA20CpauCHHR1qFDyuDbFdrrFdNto+
A6aKIQinkSRYA6bBA2uREMYATQlnW9l7INmezZ6kZ2kv0oE4rv3zpS6IaBLHRxT6rLBtKTNABeWI
S7fZCjc2CbSGtXedQt2mYfUdAsOyzmPw6C/vB2XWGcEeMpSber/GHfaW4XFLlUSgnxI6/RV0BsfZ
9EMD/Sr0aoxIErZWIbLiqirhAYd5vM/vjpTNV93oyna/hivF12I5BGPEmFpXb4Onr+BK64dLCDN4
IMxyx8hkmoZfU/dmmovCCVKDpw8i3OzPYmcVkp9Mz99QBk54j2moAsmLfRlKTID9b5ibrWkqnzMc
r7wfggTUS7/6uhiP7INNXFww5IcuFk61g0c+kfzMg1xvvdOUJMR5zVNcCc8QuUaBhOcsgHXgiyQA
TQzSe9utpLL4oIwLpZnunz3j8SPwYaVFXmnKkauDubwyMzKOLlu30Vg0gmPQ8jcdvu+nbgptkrB5
q5k6vaWpLMwx134sYiIRnN1C+tTlGpLEmvU+8krN4gR8qbzxOh/z8EECJdpsEGOjPaFvqz6lGAyx
/Ja2DLGp+Hb1spKmsugT6L6nJrK5q6Ei0PIYSjZ37BemW6HYgZIeEzoxW+dhcrRiWdheE2uFj9hB
NMebKQCqzZ/l0kwLA8sX3UM3orARNftmE+6JCKbHEBe9BfUOdAb/O8xRVwNoyJiA8WCSrPn+mzUU
qObKXjSbDAcMfGyM+8Bl0Nc8z/httiT1SPOPLeEB2c7MXvHR+ZfRXnr7oPUcaTSuloyKVyGlrhLR
cGGXPnjpnwALDmUcLr4jhrbWk78vOZe+R4qRcxWJgCQD4osKVofcfL02UqjPGVNwTVpIemERF/zQ
76YH6E7IWnWrVgaF8HS97T8YsmRDjELumle/ek2RHQ3pkpKdeMxWJI1E5cA+p7himfKMRxm1YGou
xeIUKdrb9cAymBRAArYkTkv82vkqLc8dRGE3ATiX0Y0Ra04ireTA1hsir/w6R/chiR6pXxxRZ9Vu
NbPOBgpMMEBsplmOW1Ngkuco7Hq8MHH4+WX22pLxVE1qFlydZ2mM6vKrPEPGr4jZUf0s+F+PUV3g
PSPoEmjJf+ulOxh1X+PKXNj5BuzntYYIspv2t7WCTysmG7ZPtR5MJ2tK0OxXlexthKUx8P2t98nw
LWHZteFq6Me50wl+YoHGNFwgr9iGIf3M6zX7ngaCUfUc2aGdJ3uItY2Ui3XI0IenKhjmvgUe89wu
wDWcCAoZlAzQMOYKRByDxgMgmcI8HlXVs7AIBm8EeGTwXLl8ENznmMpvBzWEPPQPpHSB3z/bCKan
+J0fiG0QTa9cI9HjY/GbjCQhtMSTYjCI016aWdkYVxtukOqnVB7LPHeKELg1CPxphcUOWFLWWx6m
PmiFkkK5Gra9T9D97BWS4OYi3vyjZEju+70zd7qMDqyIufgwN5GXlQ/U/pKdDmx0694xAlZF0fF4
VBTGTBdOI2B5KpTJu1gI22WGTelXGDXP2lAdlfGonc2JKyjH4tpiEUoy+Ft4TGJFoMjfc5J7q6GZ
0I4YIx+PH30J3pCWEQoBcgKdqCHZAOlVqoCzWhz+pxDKWJPoo5MjFab86wwdGVSDyZz0cY6XkUvn
Qp58pFRWbPnlLIvCWHirJYNLaZ8XQbOpvrNiVa37eTYSs/joNDL6FC/reqXdWkPzPVMR+OGvel9U
mEhCXpnIlrswrCamKNbvjlGp1W7LsBnGozfjbYlymGyMY6unokGkLWvvfKqM/6AENrO9mFrHMeVO
H2vQRPvZE7kX+3Vp52FuaWDEVxkGTyKEgfju+wtTQU/KH1y6YQQvRdinBigoK0JFouFtfe+gKBJy
82GMT1+Mc0boWpFy6KqmKoxB4UGzZWQSYOyw+DDEoSzCBJ1o3Ih5RA7EX7Gy3bUyCaDzs8LtP591
Hq35yVTWIFjlSLIeTCUvSi+eSrug2y6Un9M4/HQBWJuqCkDjGG9M1lbWwe2Rq5T4pZIedqoB5VD+
cAXdqO/kibmYR3Dmhi5CQXKDzgOsLu3h2tbGWcsoFpr2maWHEDs8C95y9tjNnqpjEHOP9kO5dhbk
DLMJvM78CzEMsaWHlY4sWdZgjJgtijBnfqAb6D8G3S6nLAUg6wsYaquF3G3yXD1+X/nmZLw4zvut
BbgwrD1fInNA5txngK5lEahFH3yp9j915szV+qMms4HLX2BgwEPOBXugDdMtxv4YZXq70RM2zYS8
f2dmadRcEvJYwAjMSUd93rPFAAhr+grB55Sv19l6m3p+mZjfBzlOQaWL36Q5PMi9D7slhKRd3e2B
d8b7f8gOQwum/rnllM3nJ6pQHBvfR+EYvYm+38eOiBk8w/0SLvlaz7wjh4iPqLSu0WOZmMhdmnyQ
iwlsmSydQ02orIeswPMm5EaVkYlo40Fmu9IpiVl2JlT4UWSF+cEnk1ZDw7NrCZHDHJBulsSAg5/G
xwqW7cypqI46gDnZLJErCVoYCnFmOObgVZDRa7BH+6uPKBLKua55uNM5F+TEDz9mwlracc+yg/Ul
qQifPiwob7Z27un+/GnF/FhXf5oapkF1Mzohr70KctxXxO+IgmPJGGtyomi0rxT4dkgr2ASzYRIz
ettSCmjKRkhJbAvvV1bcJAgwnj9EMrRM9tADBq71lcie5Xw7GHqVQbbNAcdYoRTbF4odBRZADLeu
YHqZm4RLUC1NfptTEVUsHj4hn3+7LZRl+D3hmttV/MlqKI5leN1hPU/EL7wFSwI1I1Y70AkUxuX+
KC++k5+WddStEd6wmn/U0A4aoOWPhSnHRfrTrmAsvxGqqWRUXkVYen+fJsPBTpehwxbieMMKMrmx
JACnrIQKu2pvJAx1NCTYqo2GuhdrVLAnwfG5UJbTgOfMlYp1RoStnjKys0NS0VbizR5vB9o18aVc
3ncocHtDsUaL4PVlgCNgAtFznOOfzcOg9LvNoXdkgXmsx7qHpSFYmcQ02RuvZBatg+7SBfj+BtBw
1wB2htC7eLGinfIhJmg7xAmSbl91/lvAsxK84oNrNHt20ghRDsgn+gMkvQOANj3KJe0xkXXwkC5i
bqyo2pNrlbtTQcrfKrDv2NcTb9ahl9HeDQaGajeFJkBZbUPJp/HhjeQqYg+om/Ew1PvNsxsxR1At
ioOiFRq0nObja1IzzRd3x1HU7h1jxkhfOnZEy3KVSWuCvH2DCBRcivY2en9+yV9fzhCFr0HGEU4v
FciXoFh+hpsqa1ook4Gv/e7G7YFCQHNNdhf4/mrxS0RLTvHPHt+B6cwxGr+8FOTlGkCGGFOqsZCS
Wy5oWf/S3r7qAaPkycCOC0n1cAxB/YVXnzIPikfG0LgNJBj+p8C/Dw8TlmvGfSetDnA/hPm/D7X0
goJK9n1I6LFV7LYg8bCSknHZgDw0YHg/SvzQC8yTjXHjaKa9Orezs20ElrCPc8rnhtWNlDTLbLJ0
I44pg3GBtW5Cgmi9MfE8Xf6OMei/l5osVF5OHX7ib4AHzWTsvmYjFiXgZKfp4KodoegF+bMMZvfA
TakYnGyobdKZNTjsNSMhvDZtt34bvlmkzW48VY/FsdDcyPngW5soMMqmAwjlmbnFQQ6zv1N89n7w
21tdL85w0Whh1hW92b/W1pklv0OD0flv/yCe+khDxFOltgYzZgGCkeBylmrIUYciRNnPbfly1LY1
qoCNMHF8oTppvB4DIFTUROqLnFQ2LMAWNZRwd2MPiYsq7Rm0MJlk8KJlJehvtGaovCD8vbQMSFtG
CZY+E2pEm3XJ698nnSq/EgQg+PgbJME7F0IKUCDPPflhPuVomme1un0S8vQ3DkpQekDEPMRPui4/
NlHTjN/xxK3SfH/xn+6TSnJreuqkNfqvmJoALO5WPcw8v5DL10of5e5sgslwd8iajBmG5z4I90nY
d2Gnfdqw+HuJ0/x5gDx4OjKR42G3k8l2XTib92Qyxm3ZEHsM6X/9FLdly2ja2A5ZZ4+vlAROzmh2
j4ahk6ZswxSvsovylkR4gPF05wUpGLvGLAU/AS3Hm/dJx0BADeQqIizVBJyUFXFql1JbbO7o7HxM
LxDlsy8eokffD4zUuFUbmhYt5GiCFQt1iiIh1W4og0VK5JN6J0U18PoC7VwMmzyqjZEoY43oeZ0w
Grsm9wG83t8A4UEDdOGxJIxg4iFKX9VEJFFF5KmWzG76cuJ+0yzpNkP60l7MMV4GcUKWKundFNX2
P+dYOUnkeWrgBvjyoMY3LFDoIRFljVfkJvSbwzIPLV4wmR29x4Ejw6ZiF8Hez+57sEIX5cT2b0at
BpiMhm5I/BFoD0KHxj5tLRjiig2pTBgHjiZe9f9xMzyDQ7ifopDPLVwVwd7sOZuklE746l7lcaM2
diH9iVm9sZX1Sr/tbZu8qsU1lwmsWyambjhDQRFdGqWmvTIWT5T+adfLLAagdws7n63ldx/WWoSD
xdP/s/27mQiZn+B+8h+TKNJpF2qxekuzwFgdgFK4/ZOZkrqEMV/WaJotg+RSThqZqjvdneSGAnHR
v9VW+s3KMKUq5Yo30iPqgB/2iwLom8L0K6Psw2MtxVwqrZh4uWkEquVLF5BZwdt/RPI2cZL+HHRm
1A0l8vbVytsM6L8yQGwHR7GB86FCrJ3T6Ock0OvhHsawBU9JsTMIyacpEJBWEL2l3dH1VbWmSKw3
o3q/nEqJrn7qkggogTLaXwDqI51mTmxvM8qhzcv23Tq17wfXcR1PUW7pZTItPFlptjCUnRe0QF3X
X/FOcPTR1ccoLQmXmdoq85hqNR3xUHe87klrBfDyPsTayYUIlZcn9qv4YS+QYKw+F1yD7Kd1V1rb
AUA7rrYa2gSMxu2gxe3rp94U4Q4muEFUsw51Nh1KyI880UEOIzAMCFpyWZUyiSzegVgepTr+wvHj
BN9upSJPEIZjHtsefnee9NTlxi3uAjZ9jCbXEmMBIzuUr/vQKGc0QPfHgu9TgBn3KL98C2GxhJfk
ULBkh5fGzK1udAB+NkMBPBN37t+IPLnUhD+wmQUpFs8XkvtLCWZAtpu771Pcpkxg9bV/Y6n8lPfz
8dfrf3PnK6t8RFGmYMHwFNAfZ047H5MbOPEIHCvJ3aiEHSYdWtXkniKvHVkFyP51uT2FguIqGYc9
O6DDsJ8CoFVmIJbIwhuJmw5nCZi1WD7ejD/pynKDJGNkxGrMx83ELMqqNL2vvvQBAFrIEZpDVmhd
9ZhRqGjT8h8R20d1sesUwLgHH41CGYrK5kScJMnDOLwXhwgjcFeNFIO8MuWZnOWyoghVcKLoBYNa
S4zOdQkXi8bQxsYU6dYd5Qzvpbw7R+BhjhIKMfmN7bNChPIPGqtIGQQ40Y5LuBqKcD85vq7WW7aA
ry+Fy0+VX5b8c6vd2ETvA0V1XI6yP70CAsc/oluemiiSS/cTIhSbU2UiqAQqLXMkgYuCrwsaOjBQ
ntwrMq7jzkMk30PTXWsJulKIEa8nTh4o5JBq93OdWACPGERg5zoxBtoQpWxdVuq3jMSKyN9WkZHO
f11ARp/1yCgc0hz6IJHwjJzCQXr15Pv+gunytF7bVgDdylJzCg7VYlL9uJnA0EoDZln7XoCE4+8Q
2XwYL15qylh7yBzzOcURt0jjzbtW/RQ8lZr7F1ZeYpYeMCw+vvS3BPebNBKRyr1v/l9P6wMu8JMr
+zEEmyj5MjdwM+w7+E2atQUVxhuACMp9MX3tWy4CNHk9N7wGElfCc+XLKpBRoCMpQ1n7TO02WqMB
UFqxU+LeApk7gFDgDbv4qEOxIN5COS8CT/xoSk+0XXPd93NQo4WR8HpJDC4afGJIaUtHPu+yV1ba
DKvQuxalAp3xDDGTYSfOMMgSA7OuBr1uyYrrhWoDq3KBxaOf0fGVwGSVy1wB9t6o2Ahwkughny3h
b1JZYQ+KuTaKGUJb2WmcFGvsMGz61f1G/Y0W54CLum3dPprBMh9t+jmemIYJXxFFyqvfnoX6qvoG
99kmW9iRR7E8lsNNiAt8+J9G3lNaAnuxItfjvdL/xkbXrAzIUDQVLY00OX99hvaIWAEJSX82pxXg
N2IJBv6rDh3b6hGw4QCoXjqiGF9YmJMtl/cV2miteDdsRbfhIDFIKy4Q/eg9VNbRrFuuu6URRx7q
OyTWk7iYrAHSAxeXYbL3UnEM5tpLo6QgLpmGWTKOcDpPpDmuoVi4wpiaYJeSYBz48c5lzBRHXhZ0
CJZIt+oi7dzC/WwnPlvGmWx7FYQwVWa7inIeF52go+qXFEmTOci0x/1cCYoTwcWyUFg+QcSYy8I4
lIuN8+0E1JY+G2onhdScMP96BqIL9+TYrZEYX6D2x/t6RN3xWXtDy9jodDmaaVrCu9BILqghMX3E
ltGrWl8A7v4IZQTheAnxwEYpGhBa/xNQeY33u6okvuLRDEZ7JRCEgsAER/Efz0omUN9zrpeB9Zay
0bYQ+3t9nmLqD846KJsQpGXtFcuaG1QiDge5E5TkrGls2fFGHYSHhs1+8yz0PrBvzhjPms0p7ofR
e1FP3Y/ddNHf4rcG7BFOc0HfcISXg1n+YQWCdWgu1d090M1W231c9B90oNa4QlkumXTwvyyzAvTr
jkK/sAJRN6gO9KfF1MVvKsRoQMrLmJfjATBjdWUUQ8v/xhMy+FwR6hZlN4g0xGwKTrYkOWsmruWG
9abUG1CV/bhestAgOQU3NTjRC6CwiY8bmeQUVrR0C5Xq8TlQJRP/KOh7eB6opjVFGbbbjIKU/ZB+
LhmPYRkn3Yp+1uzaO1TnQ9lx/MGvB8ZCKKmsf0FPPptrC9ROhr1mpP6iHH/TtO6foZuMt8Lhirk4
su/Mgbo98EAkwHP1fX+OCR4SviTER19BzZSkSMkTnPwcoBC70dmphBFgLJfw4hncW4Ue9be8pWGT
0o7wNc3ihl5iuqXMRtvWpocHqVWdhpYkzHW4XT7lugT5W+bSR6q8l6Js6lBCUpQsQhaLyR0YlRKZ
mOejH83TszS6au6JjFAvuWwK4yPCsQKfL+4LwCDvHn6ByNVyNPJ4g8IQiS0od0hxReGO2oDP4MIq
kR7XW8P9Q5JohvGI93eNYWGRSakpXKBQD0D8upNbiGbOkgAVtTxQpxRnDfTyG1ql4fOmK6WABApq
XLMl63wNmvJISJMsYBEy/SGbP6cNzFeIMPdDQ6Xpt1Gfmv38KNRw5ePs8wO1B/ZU6UZEQZov3wu1
vOhNP4X8Tuy1P5lOWi7Fx4mK5pZ7gn+5Ivub84ska99zmN0ZtaPMJCQMI6FhOSxdyRmGHQrRSe5I
fHlgFppNg6RDfyEdN/uxlysrFQwMYiChFA+/zyfO4SCyhCuRoQDpysVys1HhLq+L1pFTpGe8QPRS
c0S4DwpgnkGmVEW69uEvwM2U5v966yR0jGHQUTDHD5Ge7thz+es0RiswzVjHSjW6/JmCJ3GJtvg9
mxxOvuimKnE6nJB1gbODX3YoG7LXd1G5d7dKL9veXD78mn13R91/q39qYqp2s/iW1W9nqVG7zHTP
NhO70vsJvixm+1yGxAHqxV9vza4RxrM0afNcw2WMNhIKKupjpoIdVYDSEouLXoZmO2TcD1wPDqDn
5m5w7VNbSYGcSppBukjiFWzOSUnyMgefldXoRGI115F9CZIftz0LiQuMVJ9nc38YBMJYPwAq+S2R
aLjNdpN2fJb68biPLpQ95TgabL/SSc/OIYL7ag2omAP0MeHK9a/CclqMG38g3CxTrNZAEyl/cknN
rN7RU7JTFNSSzHeSbG858qVTz55I9gM5fs9nG9cxYCwMaVYeXRwng8Mdmo0pWwGCeZGgnQsSznvi
g83u1OzywENNH1F+wzv91VY3fYOwi+Ccq2AcEAVVPJdfdo8ZRjL7ozytRn7lNn6rh97UCLt+2H9u
9iwDQLGu1KqTnpqUHy49/JORgbSMFW8P9DOxU5ycU7jVlAbz7vPYMZgJtLnIvt0PvtFyVCTv5XL2
wCBIqbF1deg2bssi8Iy6p+REdLx0on2+i9EnF6fkwn8eIjNwCQb60VJwJQLqCq83pFqIZ1uXy9Wy
tt3YGRPGGMjzqDtgzS7sIXP5M2qMGWWFJ9fHbrv8PGtn6PZOIO5yFLnNU0cMAyn56RbIJqdsv/pp
YWo41l3688QY98ae2Bh+3q/3xF9WWWm9G4yqCdMmWvWwKe/fKAltQBS76hnCRigEA2Yg9XJToAFS
+TqMSxhp14tE+Aow2Wzm5qsLgoi9l2xNrCbFZri3YR/M6/U+nzakrG6honWcK614blKxOX9bC2Ou
/3QdvbAFDv8dkI5NIX+dL9t9qLkPoe51+4SkYWtlIVW2ntUcTbtPUyu0oKgojaSecUCbMpfgTZLu
XxV2wV443rF3g9LyI9vxo9YA29pMlpCztLpB3AXXxcyFSSvPQkEJagkWeM81gDVS3xzbmFpAV541
cdVltT7EEb6bKAUbj2qM+4gC3nmQMx0+EPKt4NYP3JwhFisKJW77XdZmNNnfxnUmHv6YxpvjqETy
AsUl3QrJO/AiNOAczjKT3ma55OchBawIxnltfWrxq1wHT28oi1mwzaf5SWd1j3pCfNLymbw/33/B
+xNiawWzlNbc/1BOtfL9FOE7y8Jlz1HyGx73GiUtY7H6POyc3cUTaCZS2umWgkJNORkA2uTvkd7S
jDrgaxx1G1oSZxwLcISjjUu8Yq2rxlLRvdzd83efLP3S7Dx3thBLXcukYqjwhMkYfk6k4FRtOZD4
BFiQKjth++Jf7EuJZbiX5EEDRXnMMa5YvDGViSXJGduEdNhG/oDQubhx5UxT1lce6l/z51p4oJtI
onMswYzdyFHc7KnRsbfEgX2Mvl/kHDjK+rD0FTMtEch38loD8Tb6Qs1s/PmodbX1sqnI7MlUshXB
GHcW92msai3Hr2hcGSxtC+m3pe6cRR+bJSWGCYZhJs4x7y1e2kXmz+qI6usksut7XJaKSDx6UAgM
eMYK6MG1SoKFSaSH14VcMlfjG/U8mz3iK9zHMkPbrLIylsGeFEsdT17LFDU+2Tx+UEncZ6pgnlq/
+U7T2F94qnoffXbdyUazro0KjMEorUdQVfkf3jpxtf+5SpJRx1+a1RKLveuy1kd87n945vBeiLQC
gOSXEKxzvLy0485cI7oOUXGgF1IIuafAtG/rs8MJyh1djYpn3lyaQvJ3jq/u61ckn2FEWR9pyDlE
wI86VTl0rF2AEM5qA0N5DPJQL5MEhZMD/M2gFo0Z2EfNOzv/xtiZNqm1n3YHTvcPC18XreeFGzB1
catDsC98Wn/RLVSL95jTkn7dS6rw4tfSYKpPwmgY5kCGfBmS8qhMiDSt1ZzAr0Ms+1BWdt+hvupH
lBrvQlM5IqoQKmzjHkg5CebpipNToyQl1jxDS9dOM3KzAo2PNyntrdrXbJFz+mLbjXz9mhCIfbSa
yaUBniocMUvj+4lNbljEmnLqWBQxWSgB3KUPpagyXso4Mk2sH/Nb729ePMqPjTLfdIPwXpeI5XPe
FeBeEUOnCzdpkQdk+PcnhQHskZu0q4ifn5XSF1GlF/sdYR0LK1mCyVYcXp/LlBE5sHFdNQlAxb0w
KfwC3RQXs2EKzzCZ4pvgxwkmQCb/HOl1eA/iPJ6Vs4XhWi/HsvLafezr7hguxcmLZuv+rxHqThK5
uCnJXZkfI4QbtE4xbnAkYkqsGd4jJtLvrDu3rN4AXi5UDwCBJpRJwvLvEfyVtMqFK74gaTYMX4pE
8acMM3pecnxbtutnANNG7vLIjMRWY0JW4O+VJ/31Hx70Y28rCr10C+4dYTTyr6AuCJkdpDMG0aun
TOXJk9C51m9QyzZ5/3mk2qGEPgChjCEVL5OUQFffyhqig0mfuaHuI9cevHPLAwgBplFyte//keUR
0GTFaDvb0Rxo+Z/27O1A03WV6SFtHf4yNI8tsj2FcIZN+e9hlmiikWvz7mBLSWId5ATldBLmRetK
jpiSQV/ooP0LlslI6HOLUuRbcmoPKOzV1jB+s93Ea/ESueXWMKPonxyyJpe2wntAFfwo6n1HAE68
2aU+raFEAr9uUQ4g7UK9apfp83AfgubEAiYlBL3FmdtmJnNttD9F/L6PrpmB9lelSugGewR3mAWB
tmMdDsnCZy9PoG1M+dnG9f8up3cSYwAoddp5sn6bj9ujnORfvMowBZYuE0ZMd9xTNk9IZCz0CIDl
pRmu3v6uS/Gi+8LPM7k2kNuePuvRSqLyH+xxPyA7XU6eSuVVEnKp/795XyGZmWNHnUewihuvRE/C
oAySwXmQ4KkEAbg7vWb1NxbVI5Tdmq1+8RmatZE86V4D8b9Jp+1x+jBMeOYw+X6Z5mFKTx3/f7RJ
Cj9vR3EEKek62TkyYJDOCtvGjpcqgClMXTMUxddlomr4g2bTyqVksD6W4sSi2sK3oYD6PA6DxbwK
IJCzfSHdx5sioQDrE4Io74JF/ZxSqkB/e5NxQxkGYvqpjzLtHMy0VYcESqSNI7hJblUaIWgWWc4D
K1N82cfgJUe8i3DBnnNTSQCc8CEONosNTsdg1mtf5Suatxs6fSfFXNmnB6Hz6h3jB4r9tiBYOQol
qoY05QifzsHvoopDm/p+r409ffBzp2KcPhHB6zwaXSLdCnrZmB4rocCYnG+28bipJoZi30SnT5/g
pXTYAyqZwVsycI57yvpk7V1vVpqJRi9pxsTZQH2XX/F2MsdHV2aO37pNknTx8w8H37h5/6hkP02I
JXFfUDe/QsyKkgOMS7SujsMeQY6jEbtNdpjoUy3J+BNuZmgxPyB894WOpzpPORFfELM+UVKyYsVr
slIgG05Rd1M08jjaqw5gRvp6sSegWsQGIv92XFVClgroopDxIlkr7XjEQMg5ziMfOO8IOtfGmp4n
wXshYpMQ0Meh2pN3cFCLmWDdyMlwPiBADLd1xknhc404v3uuo4HK1iIVKtLmS1T7Hrq0oVr8F8Fp
N66kmWNwIiybqKvRqVQEpkI+wDvX/Kmm9B9+85NeZT3LoGIVf9CYC+DeXTRa3hVxdKOGhbPDd0Dx
NRvqLhE5+j3rfjGlShcC5qOmSV5Rq6uTuaufkdbp9rgjdAweQEJOqTwzxgeK1rbzt/02lYkqXIBM
WfABGZ6JkdEsmFx2/NVGdNgkNY+G8DfK0gZVUg5V0cNgFsIDPBEDVZAMf+GLYVuW61BhWt1QBqmQ
EHbezAoGOCi4rPsWGtgQU8k93HrDidHxmED2jVeJICn4NJJuY1pw7C3d6B1T6iOqEUu6DPmv8rS+
ba6mylPl5xOBgJYRpEkvlrYkgaWlOw4PtfyTXoomtN10yH3EFXjG2mglYv1G9ad7qEaW0Q3O5qXX
9lWeA1xa5366rvbgcQrrMqlMarRuOrRJZsTwJVTHFf3URs0gj8LgLfSSH1kbEAqsTn0LL2OF29au
D7K8yMSu/2q+jyTI4dRflTvHMAB3BNNLwZO7SMTdxB4LPSU5/SZFpP3zAyuJG6jGPICRFRukkmsr
//H60fYCrCGPMf9wuw8u0TVX4lNyaMY7Cr1qIpDjVUjOOOWKURiClb+mWIYOBdkNIiEHbdZ4Gx9T
rUL2lj08rGijxE0BYcAG5Xc/Ah+3AyDKUEt4nFlvk1IL1xhsqYx0m/XlaAZlNs6kVAtqGazFWG1d
1KKsD8sG4Y0DOpkXrL4Ju/xXXPz0f4XWG/B3h04KodV/KKuq175Cr7j5vKGC3Dd1RBwP/+bWIgoR
io3Guje6h4tyO0+GTyah2bRAmnKKlU8E8tSrhFViKaDR5oSHHLCiQJ8Jlm4hEb/OC7I4YalbwOEE
4eO7yVGIzQ0RYjCn6aaqDk/IbxaF+Xjp9qWumJJqvmjb4mWBZh7mqD8cDEc9P3niTLGsyKKKZ5pL
Rnhy951h4UHGa4elXBTsiCtj6g5zfOWp9czSUsSB7khxkTpkZVQ2Yi74AZJqfH2hY8oYDyLiMP2w
IvvHUoVD77UbgeHwpxuvJfs89ZH07wKVz1MVcOc7gekC/lvjMi3oaK/H2iJYuz4NwCvN5avE7ufX
hJnaVPogySDgvnEfFK9hBcxD0wEW06c75I40zBvP+89kx95LA1tiy6F0iHWzToUxMl+saqxmcbWT
PlURg8G3thZ1F+jUSDygXFjvr15cbLE1TdeUnwoTYJFYGPclVPDl4tv25t2YKBrU3w0CSIPsUC5K
MACaeIwDPGG2ZY+LOwB1V79zoTzKTsrOV9rSHgVtOhBbAhoOancCxs/k2uI7FCksWaR8P2/fruPj
hqXbbIgZh8Yo276Q9ko9+QxiucMhvZZhyLrWfxcFdXjFCiUWTU3fC0bGsR2mTAvyAR2B49SCFnJh
e0Cpv7376fxR3vNL7RvB/5tDc3TYkDheG47wRLT3UvpqsPXFflGiCtrKocTNOxHS4D0AwlZVW/fD
joOxlEo5SC2WRQFqYB2MzXiUXeIrxNsLtzIQcnA4Sbqc0TqZ8M35JxCXRnS2DvW257Dp2nM2uaTC
qDmOLQf9e/1h/avvxZYsxn7pHVNcMr6A1roRDBjnwFa6LtAP4y5cbIdCDSUbtiC8tnGpPXTaX99L
VLRPgJC4itJkIBdhmflfBsAItBllfC2BszBHO2o+Np1ui3p42kN13K8y0lSgkbGd5DBe6jm+QLw2
fefqkxd73Pls3jnf6/N1KOBUA6glyiM7TPbPqiPI7ma1xWJwLlAQgBPki9g2yrzaYGknUS1mMt7W
XaH3hJ7T/2axNteUIOGSVB664s1/+JoK6sbufdRaklDwg39AyRJJZYtyL9uRlfEZMscRMnGsm81I
2WINDKEd8IsLvgxjn4/gUKxco9f/8vPTcQV0abM2I44U5PXCMSopYRzkgeF6EYPDrbl3V3hFYuDS
Ju/aEEWhB5RavdxgkjD3inQ6sbZ9u8ryuKigIi+CiWbTGzNIyzu70UWbiafvnDonPlk0GZmxOMZC
wf5EjY1uo7hbXthQnZTjFWOUpwVnF/VbXp/lTqoczBd3h+UsQ+7c9vTdyDUDyS7g+giZoYqGFYxI
XuqCA4slKEQHPG04GuH7c11FI/x8EyTAVONix4eRMxU3BHQZ0yM2bLcpwcwVk8P66/KbcdIZAnP/
q3jI4hjlANWM7uBam3lMljIsDKd+a5NY8b5VmcY6Ydl0sDO1vx0WtvLXUqBgvwyKtMtHPj5guibX
508ew8A8cIERIm+vhWdToT0kb3g/RV6A00JnjJjhUgC4ygoLZbfQKoj3alCcxGJs6SeZFKcS8oeQ
IJkN/A7sNITOQ1XDVzI/T6MlqGz0BBdR+177BwdeUtI2gb0nA/MvlcE0jrbRX0P+30cGCgqnsont
hMQl8kEq35LsUqsMYdtBN/DeTkwH5hcwX8u2JKL9sf6MrTrayPoDLymvi5EHxK4rnXZr4MX0ie9d
TMrZ5YixbI/qEz7EE+l+ZyHFSyc425NseZEVjXBFafWaH9BDN2VGXexDNTRxvha7GBenOsYf9lc/
FIv1coVLoIZHal9BuIZHe1VnYZgk0Xj5RCVnLZ6evEi/A/uvI1nFDE5HHpTgzii+ieDcsK36xKXU
AlmN72v4+1AeNF6DXWXdFb0fqVCqboG+0CJiDqRxQ2L5EOvbuWR8vP0HaY1f7qfcl1H1GllbjQ8L
nHjZVOiNQfk0uoqEFL4eY3NhT9LmAONrT+kosqlhWvA8thXggcDGG39NyfdzSaCxuHocBHHVdksS
efB270zmnxiKN/ZG+bLQUaIIJOZ8cbtYxrD6jf8pwoJCgnJtCHGs/qiYwE1VMmCC9lAUSt2ni12e
3FvpUJxt6TnLWOA8b61L64gVPq0ROd5Tu6o0ztpnBE2HXIoliqqS2cFZ4R/jtu5zjTakCrnnPd0N
fll8NCRmHqG04jsNjzHPHlU2CfYB+QqPbn9PVL+avnUfPA2q/2klDquSmWr2dMy96CL56DFcsQlS
UmEhUCMv5dH6Y98BekZuPwd6/Obb1Z9b02v4oAsmfI96yMIsMZm+PdLw/cFkEqzhyNARtNiwkWX4
KifW+ZzuEu/AX4ERM/ObTn2i38iatu4KluLyz600T74d0uY2e4R4zAHJRVJgJUzxNJZBMhAeGydV
02C0LTsgG9XqtaoHKyPfFMdL7U0U5DnJq9o0JvjgbbKJBuGdvOyDujeZc5uGaqk7RiD3pqEVgr/o
3rKKInZAA75R53IAPK7UGTWXEzpzsWesJRfU/Pv8dYMj63rv5z3KvRjEeBdwpKxkeXMFjLpQOw/Z
zoUJc4aOuFly/PdSztaXpHQG0CiQiECs6VuomyG1MeaUOU/yxZ44hETWSmsPW/wrIGfDcF2mEifZ
m4/gj24hgHVpecLUyDoMZ2mo78PXRg57UR1Hue4rgLLa0wn4/TwIwQaMWN6iwNtzKUcqPgbuscBv
nKfWZexnjHfibyQBMaSZ+3lCje2/hIxrXlWjjlix5qtet9onk5ZX246Cdp6gdYYdbWf9u3c8hywd
u/Sas6r9IpAIcsDbb+WDCjmzaNVPWY8pcQJETKj3fNzppKxOKGTC/kGmRDwCfQb4gkCXt6nFCWT3
mpwI9bx3uflOlm625UaeD+MvNNkLu9TR1nVa+D62NDyKebK0jjpa68p0/vsS5Zcb/3JTP3vMaElD
KBjCrPb6TDo46BCTpak7F77avaFS+L2I+piYbG6Y8mes7kw1i1VbenkddwllriR5RV9FG45bSnNR
/HA3bjE2bXddbjn9du4AbS/FoqHCmsFTTV/UEsmPQnfOZA3PTqiiEOkd7VqVr3q5zcGQL0IcPSWQ
f10KiHQW+6pfP6xBaqEdxaY0SFD8CcKiIPCNy4Ga9tD9Mdou4lpYX6wxQPaciStVIt8bMU4pyFtA
xcMlNPeo/E8xoG20tc9uJD5TFF2C3oMMyDoW8/Uso2KmDGdgifOKLXXZitL/26GNYlWEc+ZYSv42
5uxGnJ9JSwDi/JW57p+wear9cqLNxH6PhnA0EkdKculXSyqnG211IDwSbceH9JCtDG6SksbzUTM1
7U8e2I3NV/M4EzPl90/RaF+o9LBeHTkdO/BI5E7ShR/0AEOX8qzdDhVKprImfcIjm8E0phvYBt6x
+ZGi3ylcQkeZ7A0iMcdF13UQSLiCwIamfY4P1bprdHhVhLh1UA01fa5ZBo9j4VfmFJ8DqLzzW4fA
hb0DmNYeLc0FFPfh2QD8cRThL6p+Kxfy/YpGjBKX10h6f9gTa5dsZsQvhsdu+e0xbu3KXfvkfjnk
yx6swUqFqJ61fiybO8+nFgMskV1wW/lSyF1P2UxsVz3LwncMh48EB2hmQk0LCzB+Dd8kxHexIUYt
zMgxZjcqTem6h9FC1zElZYGwLPaeg/Orjmm2l8zxso6xHHJuxDLgS8D8KViM/PJWJIbOt2Ak+UMW
OUPQin/h7zGOZUNm56RHXR1c2mEQ1aHPdfDJqRDQo8qy5PpCisRJ78+MZkN9Gu/veuiV0AgmpEFq
7UGH+BmPLuYCn5Skyq/QPcFuwAXDNvLvnZGyR0gSqMquKOJkxdUIoxMHVHd/cj5E2UgKk+bkhWOa
B6znrJD9nJQYrA/AyAI+gNkZt29NRx4LtnaDp1ELecUhyH6W9IObuDog4Ml16PoN4cN405Ro0yKt
JhhaXB6AiwfMvcQJusAb0eVtcEvNg7Dl3wKx0Ycet0R8wzu5IKkngaWBipb2DtcSYNj6ElqX2a+W
cYTTrNGDNmgKrfifQ6A+t0Vu0Zam2kVpeXcTNGubFF2NszJgW/oL9tUbmryybCFbIi1tqgpnm8wd
Hl++tY5XWRwPO9wYsXgvLWp3QR72Q2L8TQXeIH47S+z/OPsXhNFSu70KfIHAnhrRsC7cR4sw2x9C
rqklElmw9YXxayuZR0eWJbEdfAhQPUOW4NaRiHNvnkdP81bmQBvyGZeW0Mpge19pC3q6R/f69uzA
VgWslV8haOVFjvoaPQPIyZXIs0dBsFwZUTvb9pNjkxo9vaPx/WzQDU34U9jljrk4JzrQQGxDkWd6
ilx66FcsiwbvaCtkkCtbzLAG15BJsVRZ5v/xnRSTpH1DZMH52wgdp6FEXTeORkd2ktXJYhSjtF/J
ZKDODONehLqvrlQ4J62S/h1ybBUinJzhZn0FaoFid9kQrEQQcdriksSKMgwkm+w/aAFq/mACt1Lh
Gd+TTRhZa3kKDff0U8MAbjwyjLX+dUAfl+ZK48MzyuRtnYTrEPdxRWLTz3TlhgGtDOhZdJO+Cqz+
ST2nyy2DiijbqPaadmteCWCVoXgwQ3WY1rqI2VxNo0GyQszs3SeXAN2IMn1K0ZwfE3G6y//nwYIA
e+lDeMzZHbm0bsMAYqZp/ygnwxtma+IocairRz3ulR2EhrHqZ1SK6Gzj5uO6hqOU3eLbxAZ6DdSk
wXw3xFp8U9k7YPNEXmd4oLLuZ9EiwtzSC7L6E+49LaioztyfL4XU0Bcv9MJ3gIAOFazLOJFnn8Db
VV1MizkCDtig4MovdqLYR+ZGmIFfldKe2GEDhGWkS0GoTT14Bs/KtS+25e++AAXCCqAzzxNSxcmk
9a1AX3ATzan75iLgfRWGV9kuyjOdaCV/ETN1DANkk8BA5Jj6ogVr02zkSdmxNT2cAN1Z5IfkN8dE
n5rGbZGcQ+uc9527vFOEmhoKmN8iVZ+5aloBoViMsgczBKzHi/OR9NgXupuxv6Tfwo1AeMyGEtIR
Xcp/SBC0rglQTplZWpdgR3U8A+gWkWB7NDJvh2dP/tEO6GoxCdlLEyvEC6xXuWd3WKgmXWor5ses
zLINWL8HXoy5jYUTUHg7bo4+MifvZOfKM0lDBGFP1tiLD2J8L9T+S7cpN0SMARd04pAZiqkB1bOR
BXCSqj6BlNpiMH0QDzDK7v+DYmGGrSO9Zm37kElnhY++kfb0nHAh/C/6wsPRWwf3L9ZyqJSkIalq
qfZK0ZSI1ROFMLABKDR9laNxZZxACElDy+lGhj/wRCU0x0NavzRlkWIQ+llZ+u5CooyMSWS2LTLb
M9KBuHVYQSlkpotVU+/DrneKBCGg5jvfLjwLcgvVKDGVdqgbs1HQB4tgNcV5nFFpyCCFOWShTZUO
1o2en34Qh+mcQUdpTdSlBjNvyM/TB/xGuv/RRDgDxRBW5MrUf/v8OeSVuE6Z13pSXQnbCBViFd1I
2tFFpTl6RSXWpgLCw/Hrj4m0+J59F3toR+tzH90xqg905zRB+1R3E+gQmOJxNllzn2NvcYZWsqgi
e2rtHrxirlxtcqCNzzE5M2NnPDymm0RNfN+pYKuDgI7Iv0M6MTZySsaD8KORHc8Vnq93BDvt2PSd
pK7vRUJbNph8hEU8K3rqC6PsExp288IbojKJhvS7fP/Cd37fhXC/6Q69VWLwZiflAexrlvZ8rP91
SaiPryEwMORTzOk15c9pcm4ViUVcY0jpk3VhwsDIAZORp/rB8PMq3i+jtdz1C2P1sG7rY+IWhe70
2uIC+IeksoGL6rwqpXUoKnin0gsrDdygaOcsrK1zc3uS3V/OQBIj5/D6RmxISuGHMBeBoac/dxry
BpeRj1DNdd9I0aTaRgpy21N2qtssYjuSQ6s3BPFrtzpWek2b/zD5LzUH0PAkdqw+CDYDeXXgtHh8
k0YZLjeUsFOnYYTLUzUHyOteFN+HsL5uIPvc037zrR3GtHPl5UVv04UxuG/ge6tNnUoUTsBTroLt
zkTZUlLDRSSZw8h0vkMKdGjxSSbaZjt1MzqRLcw+jEoRwCHqrwyyX+cbKTjqtUvrHDQAc8Flj7Tr
LcWEC1OoCQPi3puDxXjdkWZPvv302jVIUf1LN9gDhLJkAr+GXaWOqqhXEN5HEpIkVu/75f3YmbVq
klExxn0V/IobrMiCsWDpksK3eEMXHiIAbK8CsrVEn3/yad5NUVFmN9LNyib6EXiz/5NdKnNI49nn
V6EG0pd1gFaMOwDNG2om7KfvVsw7q/Jyuz/cm59JlLML7BcAsPmmDmHSSJhLEb4WtLageptu95or
sB6NcF4150Tvzmw3joRS3d66MX4yyAc/UIfgKqcD/FzIL819xkSE8reUuhnnM5M5vmf/DKEr7KQG
NOTS3SMVNkYxnEcSVvsVKsYk34SLbIOoIhvDE+4yh8MVWVYtuIRZ2x/+ZffsVDJ0Fhy6bcby8HAG
ZsFnIJpR14ENkhy+XfvrvrLBLHkR+EFppXJbe83gXI0/+eQxFOGpAQn7h2mr1MzyGqGsUM9BRM2f
4STIlJVJmL5FPXIf3uj0cvtHmgZVDKms9q1dxr60CuSPMDf5NCQzRZLv3/XpsbfhtOE6LDqCW9Sn
/kmlQhpFRpp5h6qzQY+t63HylRT1k9Ikx82e4ABuqyKeni/sqEQAW9389Jk98k80GX5Ql4dsjf/6
kFqSmVfVOBrfeigXAfJWeFb0hxojbTqeXp7Ikciwp/1cgVP8O+Q0hAfVjAHZPxDZuowvv5ZxKVAm
8M7KLyofcJy3G2b7IAa9gU4BpPn9QOrMRWGhCDBaxg+QsTzEVaFjQgKIMLjtVSSNuUPplB+nc+vK
s2kW+kRecV51G2rSs0o+BJrGkGGOjVgK14O/RMffPyXPJ7FoEMbUhvpoNfG1vlrRD112jqXASf/A
u8HWdzjyDFac6/qm1y23F3TsatKhQyT/Kc5A1pMhEi3C7OgmoeIb42KqolvaoPJd6Mc6TWY8Akm4
1WjGV45zyW/SlkqcvDz9ALUsqgQY6mit39oCn+CEtcS6d3xNvh36Qvx4DFT7jpluK5MeHbEahaba
+h4xiIH/NQeCIutaiWO3Kkr9i2w3cGbl+YnKFgendPXO3gnN8y2p0yIB2hc5XkF4R47t264dLI8K
OxK4cqrMtpnmj2R3xlDD+XDSAW6EekAqt/PQN4gobYvh/36P32JedEWjdfX5vbB0vY346Jax7FX1
B2FNKZF6J7ItRcrEADM2Aycbb9yM4jBEsXjv2vlDnZj8BzD420kdVt+kZgNcSumJPDckNc/kokZz
co1F4omTagKsqD/rSltxETuwsSuXCvwaLjjl49C6Wg32kyrYn8KS/rUr5cNl9WfMbZNKEKokTDOf
+qpEVEGczzaMGB5rbfSGv5OX0FUH6dZZa/azA+bwb32RdDRuMGaPQ46QtYhEcrIwIzPricViYNQN
97QXLML65Y0/Y8NOg/JqKXsoWcg6GdAPxHPmI1s2tmZ1oD0OKkAqS2JKe47BBRHkbWmwUM9f52tz
AGq3i197dBiB4Km/j9rAnaW6dzJimdei+TlMhmJypkpmxaw08ZcV2SU9Or6KzrJmsVvInR8hFHB8
h0DIVjhUptjwZp/GiJ4AqEAZSU7m526uliwXOfqcqrHIWE2Hwy61rZCIlDUEXuyj/HPsmjg70Mn6
oslZI9tz4rQhnesOCTeb/pJU9aGerTyDj55EMPKNT//w4zApihvsb4DKsqgPw6W6wkxqIOzTzhTp
2EQ5+EkXCH3UsRrMRpOWRF9p2NbabdXV/t58zz4v6b0FU5EfujmaqmjXpVthM87T9ktOhAbxbiI3
GbCgLzqDDf8OStiVNw/coRaJwJy24h5ns5GsAVUDJsUCLGXnt9rSxWI093EaIruUxx9I1X8jexBj
O/0OuFHLPgKYS/CvaA9itTW0AyWlreg3YK0ygd83bor7zS2y/vPGj8heguT8PuB4XfxfgNZtGhwj
cQi9LGNB7ildyoodVJ/967V/ejvpDAYp6oVCLhR5TpEUx1AMRpMdaSSqi0ZQK6EsrYG6nMyLebCn
pYUWo4rJn3J1bxQrmxDkg45aBT22dV5cgqwhJp+htAGOHi9xdOUHkUAKj9POWz8ztlyXad8uX9An
3nZjezWPlurVP/D2mn/5IWk0NvOqaX5URb1yDiT6FIMyxG0trpXOtij7vGKCeUxrnKQcSkLh/TEa
uQaclVyQWMCmu6E5F6FFd+q7Z/6oBOpM87s0GwpM1TSVSjVdag+nkYjpNNpWJFKBG9sNwwKCQcp9
ZRSyKklizkZKmErODUd69LhNKbNaHbws8YFLfUPhGAcKAWpy7//dgl6avMtTVd4qY8TntV3IuzTn
YOj3hvaqYsiyXSWeNkTtj6jeeKzCIaNVKW2I4jwX6Np9uTQ/HSMToGs30gvDohx/0PTCBQUWGQgU
cfalQ68FwbZ9uG3D6cAjNNTOToXN/LjVT78QZu4gUSCIczhAtGuQi61Qdcvny8JBfRlIpXHcJiNq
m0gUrklim8H9eOFfwuK4iO2moaalQ4vGRPxR5SQt53AnJC1616FWAJLCJUUwXincNhazc5nkrpmf
rB/d9jZng03DuZ+NwijCc8MIm5eHEYpeqFM/K/cS5LpC24qmEqJjHHb85+aAUP6JQlFTsB5295BD
+hilB69+2UPSpVT+pU9jZ76qR530LMc70X7+2oPOBxXS/4obOT0RJNFtU0Yi0cZDpIKOLXP9xPJh
shQxrgnInGKfmQeRMKZvw0as13oBRobijzKZnZYOU4RYpXtDvF5iet9CIqk10YEueGdPLIywqBkX
BphC7Yw+bAP/fz+4U3HXuyvTaiQ/7pr1b6N/tW3BrusT1pOMYkjaVUEnDEL0+bGxTMwRx4YnEuye
LCwoAwRMLU11T0lhLYRNys324HY/WjLZrpZ2iv0BnUKSy460ilhtFATwlgHmmH5eF3ibnIyqoGj1
ic7OnmwOhB70fFV0dtKHtG1vl9CVcEuvZkzB/MgRPbaXpLitH2ekZaxNxBF69LcQF00qdJRMx7En
iOAnZ9q6RYSoEfKK7JXpk25uVCD0/1MnSn8+xBGc3Vxy80LY7EAsBaZj25OakQxHfvuaVEKm4fcK
k+OgzGQcfQfy63Gb4wkLidiqLEXAAHIam956moHc724mJH3hkd8AsZCspPpSGuwHvoJAhKM3blnG
xjErG+q1zZP/HEHjspqFdYNfn2Leuf3aF34SGzB6/3NjKVt/LqgbUg+sb0+ywekfdBLbiOO1e/DW
p1LrJoMEce2NgVdOYdVt0ejinjKuzZ5DbZZp1JCsC1CExoc3LfPIo0hfY+9qEYvVZtnM4rhUbrF0
/uty8sZf2UjOxMcW+IqP3OIUC9/Mu9CKRdk/0NnHK2K3s086Tuwi/l6O9zDzXUsq7kHG9fG6JfMt
kRRWGF1qYqU/B0mrupc9a8z5wjr0qoSm1UVUNGjo+/ewDN5zAxLpOuvAyBWb3HDceAdAY8jay9Pb
0h9MtGBjI7oaxkLw94nwmL9QiAATiN0EQ8jopSV9jGzHU5ZLfy0B8XeKH2k40wXn/mGDWfgwfjrU
yRCJJS/zh69Aa7YpzRubW/xuvwGyfJf4SpJjyXsXlFm1ZmFGDp21qaYhlSgJok3S+Z4jHxX7eeEm
r0LcTbhs8OdM03VW2fI7HvfPQQRZBE19bgXIsRJB2nzB+WaAriBsMVnR2IiBu2hlsh9vxo77jwnW
8CqlmlIAdw4mDt+uDvmIGEl32rWh17k1yusU0j3lH0Dqx+0aRoYAh730/JXkJ3N9PgC234EmWlsv
ihuiy68ou6MqZWTepTmyRf/XxvUHQRmz5v/vrwRz5IYlc2Iix16TctLDGnEz9RIi/sMDn3aIi3DW
Vuon9gPURSZCfMQl8jyROXMboJ472516GLdhH7IZWFZqhkT3gCf2xbY/0Kxev0xBnoLrOHVZKZcN
wr6Vq95ccB/dFQXyNSnIKuil8ZtEkoWNrXBSU7rI379EKFXh4dWI+3RIlMKNxTj/hPSY1oaaIn+u
g/jQekSa7Zkae+sWt838WOgQR/GIZjxD+VinBH+nCzb+RWWqc0J7Dg4qjnSzIkdQCneLMwW0e9Zn
FPIG9f6mtE3/ejmhnjWlhxQh5tmJ0tvcUwd58/jmph9TwnXmQKuQHcixtckzP7jqHy8evX+QaG6z
QVu+OKClsHI10WVwvIiuxjLSdMBi4gCQAg1KIlkrVAhK2Y4s4KuWLbk1/t/o/7wbimizX1zvKE+y
B7I5dsrZrJVlTNGVXkjk19cjhmy2ZVrSONZ1kAi2cejisGpuIqP9NHdbZhtSfShZlVO8tEUCyD7T
IkDYpEtttARypvHK3B0HinYnsenTfJJpCCo6uZHpIyiNpFKk0FCuEg2iV39Zh6mtqf72H4eR0VYB
i9xPEolYq0k7hSDPpMTwmaY/jOzEyLY6Z5UwEqReI0SRYuGOMpfhtfPnRHyxvEA1qxptUp7YAVfg
Q9imzrWIk2gRLWu6/stmxGw2C3JczhG3gtVc3a7+jSjN3HecSv5uFuuhA42Wb6bLxFSckormaEZh
kqk08saELjh1R1QiNg1VAPAzVVqpz8uhaJr7vyxHDp+pE/5a5oCmrtzvxiGYrXBR5nctVSNxqTQB
Ny2tuj5YIHmGDSzqsNNdkc3bIfpp+UEzVKLxbDm8s99pH6kzw+1oTMto3IJL27RNy+oRx6htGxHz
limUm9+lxqDBfTPYnNL28mDuOPd7Y9dqUZb2ZCcfL6X6aKT1FZRvyJi3LK/W7ByIvoVPBFVgzroU
x08raIWOcJlCDZXe6eI7rxK4PeNllvLagATNLpxhiynau4nVf4n0HTs9uq3FuE13WUGAK7goTyDQ
cNtPtkPTX73i3FIyJUqCee3oonF8J8Y2z2j7gH01NgshlbDwMM809qdwN1/sg7857wBTsSlhxsT9
+C7C7f5X6AB+mEjV+q7Guw8LASJSKSyAwNyvfykumN9o1nMdCTXKtJacPLGC7h9pcG5MebsovUFX
FNi1jjCxh5Z9KX5QdctRcM1BZHYCihHwAu4rW8PlwmwxZXx6OGvYR0Z0bUdfQ79DjFE2bzcrqAHq
zdjogUcBSLjjznqnxEn3VYjjezi7NmksCfnDP3CXxLGB5pw77EUtzGYNqj2o0ksjsdQ/ve+aVmOP
Zc0EJ4U1sU22SGZmdKwkVXcQC5OsROgtphR1fEDY6g3r5lzHQLZe5IL6U0mhMPW4DbmDGJdKEO3E
Zo7AzeoN4QOA6vVZdgraFLbCCtoRW5SLDh5LM4asQfMjIqXYsigJKjufDfBFzYbAIeygmZ4nWVD2
8YjbojVcYerPQNaq1UPdJwcRJF6dKOTyzTBOwvBKcgmEbSQOmx6d/FggryboyY58oJcqD1Y1/bNo
3HcofyYOyOvbcV9UBCZ3eGyRruxLv2Df6n7hKJ4lDEIvtdSe18Uuoa/hPQDe5s3cA+ShUdPS02WK
50G3I0CxJLkesvE16b5mhhfJsxTg2tyUvVLGW6f+TmRyJ5X1vgr4JnPEf2vSliJ1q0j7brnAiKEC
KqlAPjYCCfuNW1rWREKucXZQ3z7prybTHbLQOca8iHfx1Ri38HmTCZg7Tw0nCKzQPEAOtcCNsCHY
rFEm9PGhhf7YZepwhTwDx6JD/fLaObb/mH690KLD0edCzl03LKfd584UYKE7VRw1G1572BiqMNuV
26/Ic+Y9EzDJejYyDCWXkUNCEYnBj+qT1yOcknGcrBgDvaBF7/+ICpQBM2yiIbbvZomrEEojRvIk
wY/ZedDEaS/F/kiGX3GxTVPaGKRqeA9JwuKNHcJmebvTqaf1s7sb8jTR2TTN6g5yiQLPEfjRohQP
7KjFSCfiXkWYo10xaiAk8XeG8k5hCuejgjb7hTTpP5BMqZ1QWADaQk5YV8RwJiUJ82XDoiT6MA5s
RCKtkGdqYN+FQRGvMzhePqBALvuZoNsPX7TiGa/KRtpbeWy3bCdWYqClYIAy+MSWeu/Bnluqudu4
7IWweQay8GXLyeGAnZj5y3PlttAY9Oco6hq95T/XuUr/802HAV6DoElM0dT1QbOK5NXdZi3rtHx5
dAWRLI6n92fqmbfAEZX/JYA13O4r5eep8DABkmD5tPk0MGiHXI9uNmIgEPtxnAWSZW36RrOMgOpH
UsVp0Hn9c4za14znmG/+KJP0qC50BBdLIW2C32HlviMpX/rrmxqxrFUVv+zM1g6SBwhPys4a8Z8L
CoLq4T3zXzw74/RolupeJGpwe/76yl/+CdPJoxOAWx9heaNBafxyiFcwax1vu/Hneq98P9f8vRNm
REvA7Ofx0yxA2+x89ffnNoZ1ubripbbgGsi0Qz3Q/uKgqb/ARfg7kVgncfgyng4ijA16S4YfzAZp
e4isCuGLsG0AauYFss9R3at0Hr+lK9Cx5gd1eHaB9boOBjXjt1Qa2eJi2TYT44Z/ZqW8PlSYKZG9
+zHVGY/0e8le16O/fdYyAY5m+SiLTdQEmb/av6WhOY+PBc8aqui1H0qFZfq+Lth4iDOqXoLKXfJg
3VG+SgNjbv3dq2uLKIEbd1DjI829xdspRrWMWV2pgQ7XRHKvNnUJ/rbt4jGFUhRIn5yd0HmgIWNx
NzYuFYsuSCWOTglVp7NPXtYoOVHlQDEN6zkvjfIQumzrJdzmC/Dk0Ws9XH/4PTgeftcdtZ8vS/Bi
mLE8rvWq7/WEGxGc+zJyg4zzwlirdLK7t/rLhb//il4CnkRBNQD1DckUsA1f0FjoIp+RBdYjN2kz
aWBDSqoY74dUXjc6KI4WF3HfBjCpHAIuAd+BSUrgm+9eciPAz7dNq+5dCT8t4cbEVh6hhcsyW/6V
se4ut14LNm+u2HfWKyRWp6TKz7Ly8HOr5UsM7MzkgQJDlfxifaWNPGx3V6uij4ooGLNCvxKCwSVW
1AA8JjwZp+eV0vWaUdZ3KrWHTiGv077wNAKt8nwk1v1Qu4QAEeDY2LgF9Euo96qQdaNuF8L67+8M
Z+lFLAdp+dcc4BxhsicUIr6XmAnlWtFXNR5L6+lypGI9TwTglh4jyvG/mkddnNHLGUjHOZmW/glh
olCWufAZIgNZxvW+Fmuyi0g8VatwZp3fGDsSeXPdMTDbtYANSWeL4G3dEWjegiqKK47YMc1nlBN5
UCCEb5rNB6pq++DlKn0Ml4x2OPBGSWbkqJlOkd3fI5qkpSa/mVeR2ej0USHv14VrUYJTUnSjMEQk
p6xdwtWLJSay5XACnT4m+CrNlREQmvtrZ7Q06Shdvuj6UFo4M1PeFzxp3FoeYlJlVcFMeyavfyeY
F5NJC6ylWhVpkMhVTgS5KgRf5LRtGVQG5BpLnLNe3J0IIYHUadYLm6Wx/cHau5mvOC0USPOEI6AW
ciCkzKj/hVs98YcimrxmU/Rq7yOc3UPKc0T+NCPdBJh5IW855BGqlX8F94xuCJ118LFnhDU5SYr7
t2maackTC/WrOllkphql8pyAvY8Xo0btZ8Tw0tQQob2xscAvL9zpsklY5ZGBKeOmoveC3Ugk4N2C
7fwH/LwhqyEgSxsCdgW4+zgGjUY1xOijx6DAqI1Mh5fsVmYxqRf5e/RD96WFAaMIFuI3EXcigrAw
R8pTqWaSdXdBjtqHWBdtsbbtAI8jkUWFe4nbxupnpfn2NO9ooqHVFPtz+23/OblCt2OpwEBEqk9d
+uGtfu+Ph4Z3i05ZzrHNrtqkt+WHyrJ1hz0+9poLAzJZjvPpNfByMJ4B2bTuo51vsXD3KfXVVAE5
IDMnFnm5MdpefDcX1uMEprqsZzHCxi1aBmpMF6qHbuDghpu2z7rpeQoDdJcZr48qyZnj9Emk8HFn
YRre9Nil0SoMDqZvMtIDf/nKvy2g1PndZbhf+kbW1sjx5evIDK7Fnb+XloIlytuvfXbeQM7WMe49
C99N74DQfKV8dk1KorJMav5SYc0+c5JZnVD9J0njKl6fcw7deIV4R511DKDtizrHdfWA+ltuO84E
QxiGl7ZwwlZTeCXiOFco4LsAtlaqOz6zJ4SlnFqIHPc1V1BB4p2Esy44mk0g95IXmw4AphGPm5Nq
Our+H3cm0CC0v76Ak/tLmRHiWFZfz16ugOcvqZQrVVMDur7OuRHakzCDsoJBF3ZY2ZCVUslck6+H
+bS4NROUCJu4isMW44VuhS1sl61eQKB1mKzUrMHn3570iXbi93Gbi/oU/kfQGImPX09dcssCxQog
Rx7pcQDZwNs3sZQaC2FPQlJF/XKNELsE20rqNksyQdvuHCOI1OXMupQwNm62xL6r55wLdYn09oZW
bfs/goeuQ66Y0OQJ4vvHV7XXlnwEaVS4zKp8EfL5ifwogPxtpKtLZlevu03THUyGDg99jxaiw+UV
4WOY3V9yghyynfBSjVrOCmCJxXqa6EPMuj8NQdTCACU03fvUMTIu48puveE+3Nc/ia4KYYh+L+LZ
ZXwGm3aTJ72rBXQhoAk1R4xM87iGOFp2aumd669LlfzITkKT5v1yJ4QYnRrhZCZMiNhVwWR+Y8Od
bzWfak3fu+xfbuKlut5J2vSMiCIso9I9JSNc9s+SNMLorB9w5i5nGCqQ9KmnCYf/xmNxddz02fMN
ABLSXTbe0IRgz7HHCK6V1f6GhgmBs0VSg5rl48ZNYiOYkknoezKQgTi0ejZlCCJFPjXXUsqiVmNq
Gwdg0l0ZusqltQVuCbk2vOsAwRAz8wgbwOnmMfpgCPYYqX7vBitz77kHJeiFQGhvvIA2O5Ad4h56
8xUmQZtL8Si1YPanM8GhLAnLFzytlCW0BljBrO2ocT73cSnYgSJiLmGwymcjgMFnRbUn6klZ5fRm
rHtHdDTcAzqmbtCQWz3jplhcmajF1ZaIIavc41ILZ7C2QmohmIJrUmZs/DEeYUatLjt1kQY/dCNi
EJpoe/M5Yh0fITmV0XUum5WsPtpr7BBx6SrxGIi/3vUAejcOMwyO2YXA7moMAeyndHUOeMU2e654
B5jaBMuOUnqZ3S/7qQ9qbtXqUjhmhw8PYo3fO35DCSlOgDhTyh3Iw00FBC/8yeS6oGe9/HHE1nry
fUjcVcD+RrNX4wYMCPuoDUwDy07xaD/ecUqrfE5txNDNh9JA7IbJYbYklTFdg6Kmu4mcz3Ytz0bg
bNG+ZxE228d/1xE6U4QJCsOOO1PQm989r1Uw4byYO5oKV37DQcj/oWW+GfevUi9AR6yb9V93jxTP
uAAzKziceY7lzzkpA00fTq6wMQQ9l1SqlGeUJQMAsDVRRWNGFnmgOfBZUrKEulwQMlW0jWegI9ya
qtHphskv5IFYmSeLIMJa7tl/NPi858uo5J87Y1LV1eBPeGeishsnowaAiHNQRrKcj5ukFeNpXNZy
OycAY5z9rwzPvVnm8/7ezbB/MZ2aDvqh7B/8lnufL5Tokc183kWjudz4f0VmNHislJxYpi5yciT3
8tcV7WdGKu5M+Uza39hWlnDYssj93jmfhvKlV/HEk5XxVRHRnZmRjwCI2nMxPMaN2IAr9yWHSUw7
/baXqkm7PwxeT6Tct/RzyjKQHNMZrdUy1DO6Gwe1m/LXA52aK+UuWJ0BoDmcAG5m5RcFJQLOWxxq
hrK6cXjWKfKIAmcdiqDyNz34lk0OhrJ1fRMTH/qnNz0vBm5i0nIRZub5VYkmUiFAC+XWshf1st8F
E5vz7jGWZFCcmzVCnQqknRBDyLd+SteEXapEwGdv27bzyNLVw5QR1R8lQFC0e50d4TERudUmbySB
CKAerpysFDyI+alcjsiUgABPDbzXOTD+fcON9YzkRQQaO/KpECsjJlWm7bg3IMQK+FCmPswF5/tu
bA/0K6QAql50S77kwpxwHM6DbHdD3b550KhEiSK4FAKr9ADstnSWpgtTCNGjegljYzfciKc1u1TA
JS2bp3F4kTGl3pUmsn47FqyGagWJCCdTfZfpmHgT7sobmohX8AedRpYA6PVDmXGzcJOb7uQxVuiw
KJbQEOr4xBWRUOAIIzH0B886WfHrDBMPe847rTt5eOb6ov/M1RBuY2ZSJWkg+YpDNzhGNqAeTDrz
UCoz804hhbyVwoh+lz2yeEbrXFHW0oNR867FvGs+p1/f6OZPPADubP2aKq/ASE1TmJh2b84Gcd7/
XwI1YBxYYBnsa9LL1Z2sOVU1Qt0VSIy6CzeLG7HMAwYyyxYEQiDFLiwRbBjflfjlXRSkve5TOpDu
1Q1BSk/IfaScM4rYo0uanpDZXu8V3+2LLQEcipkhVpbh/3TWehahZ5eajRiaHXI9qoZDqdWJbrEC
TB0G4VIOfdjd3+pvEKTqAPIfjA6HLTXkwcTCTpi/FprDdG4eqycIc4v1bBQyFdwpiYT3aOgv1Mlz
h0nw4CXjJtOzG0IZN97dZOkp0EU7jvZR5AZNbVrY7qitHxOEsrMiLzOJljSf4pn34CowSqQMuVlL
Lm+J8ifzKopfNZLE/DgbJg6yt7PAQ68BzjRjrFK7rFRDSbpDdrpJki1OYwBtA/9m7096dgGj32Va
sD9q9KJtkA5GI3WYgf8estHIaLQmLv+IdSS/W/kPkLSos/XWR1rHTI7XBvsg8O30tLUylEuGYzFB
nSDkJ5QMfLfb75V2816uPAPA8H1WamkBKbhoOt8v6CB5nLk9KAWiK2EIzHy1m5CFOkhvXLr6vETc
bHFVBMkjSHb+7S4GhUtaSTMfkk6WPzlIhzCLTLGRt6YE7Kr99KqO6U3IDmwggcnEQ3S9V0/oRb87
8aQTWZUUg7Kr6C+LnH03iunbUbbMiZqPM+kdgaUvDJPqxeVZB216I4ObmW8ctFCp5WOUanJCkJ4e
6tBQOy4TOSK1kHVp2p7ZU1FZ5dC5WrwB0E+/wLQHNsYeP/N03fDxN3waCtn59Rjl0fVAaTCKigZc
QkRthFW36MM/d4VLoyoRESlCXKFG/epKCpsdzILegNJcU1qCdw3KG/cXq3mVbkAhgNBq+g4TLLnI
ZQpDd8OjI3aXAoUfEbNgPaW1Bx556KslrV7HK1yMIo+OKgzWJ4/Vt6GCZLZVuKdj49v0pLU3Hxx/
IT8B6Gnfyy/NpbtdS9eO23HIZStU+ECqIoASaoSGRrK4Qvi64xlV1DKJwSYKJDxNGstuRBhEjhCM
qdTlyzhnNUXn955fIzVgrJTftarJ0i+R+c3I9oGu8tvLbW5FhNsLC5kS1DXvbHUW0Pv4pPf/7cBl
ZWzR51FBHSkVlu0m583n/fcDc6Kbjlt12Hb8//fc7d9390nQ96QCz4TdQxklINoC71FuZjept3q7
ugKX6i7SW3YsyXj+dslQUnjciEuvWFV0k9tMaWdUupKq/Kiv7ew3psoGHw8SCyrOb9Doew7BBIO8
NsVAVnHmMBjfEcwMmosBKORZ/6iaUo1eZpGvsNNZ77h8fVcB0lBav1lwNzn9j3GnrbxdABWSWyyB
RgqHTSRojAqG3d3s5DeupHxF+giOaIeXMoKAxHv3+a1ckiZ2mHSZhX6X5K+nR1hwLUCeEkjM3uVy
9IQB54UQlbd5d0tDRNZQ9Xd5BnqZ0qxIhC1GETV2fC22ttBRgMWAbglHqAtvBN2Q4ouFmA8oZRpb
YJNhtXpVGDT/mo8NK8Iz6XFb58/BfxGLgecvYOK4eWlM4QMwx6cYE2LEBSP4V/XEWm+zX+kqjqV7
kU9IVZ58V37XFQbZDU5FhJ99OZqvwo/Bk2YIOSHgh4iFk6oTPsfTRkMLmSjonentwevJw9HoKBLx
On9YeNeSaeiFm5IQsIDE1j0Behsd7DyXxUO8MjPwVwQTTMmJ3YmAUxgsSGPYZE57EwGRQ2A71zgv
Tf/b5vsHjxdHlXvtIfJJ4nlIrTulsynG/jnqej6wTblTE4djn9iZD72fx9RxlZDoKNXSuYJpZ6sj
BvPIdqeszdiBNEzX3qCMs8jJHdCObTt2YYD9iCwGpJUXP9udlDRi8NVsxXBAPdclx8VpsEeH1OWd
nwhtsJdPjtmir8MlfWOahjczGZYW7v6KTs4QaUfU2q8DY9Sg7I/Q55SNeGObjxgplz+/WPqodN55
0RDdUc7RaR3QLs1EvdL9+S4G029DC9e8fivstUvgmfYNjve+89CArYIjYB6Q0OoAyhguvZv30eJR
m5sW4gULUmCohdK0iHvYDmW2ywjJN2Mc4tpQdGqQfdjvrknqBBRggibu2IGxCSPQRpbsBsfKsecz
2vKtuk2lys60XDG7YiLpg2Lo9IJamddVtkU1KoJeAp/ATGflLRudB6X/sYg97Q3LqzHzWhuf8BxS
xw6gONY8cP3TmbBPyFgHqV/ds+ouIWntfoTqu9ZvZ6jnV/qppI65q1sMDVA8O8JNB+dSJb2xBnRj
xvIoF9eJyUKzRal4FY2b5Q0EGZO16xmBq6fmC0qMc64NUMP24N0XcbkmjFwMSSp2/WpK7q9Kiy9A
xjIXLC0ig8gRwDd9wD03PwOlOszEh3Lu4hRV3UstYAe76rq3mOrTnbacJhlPLZarhYnrizBkXpDz
T+xe5+2xkRld4LQLiYQpKEXqIH7BdzkEYqJLfUuBBe6VRXMq+3bkR2W+2XBivSUO/Db6C806Pl4w
Nu0dPAPywLNsIm10Q+z2mgIwIT38UmrSdLXCvCjlxlBaTEgQTpDjxYVA09FNbP9M4u8umi0QH539
1+lOEtEm0iTK+Ou2UaI05CkYbQh3D9cp8iaRgDVVmOdhOZTWtzlWJaB1qHjFXygWQl1rJhcP+vaF
PBEM1b2HUOgR8pUMYKEZ7aX22imGy3tD5MshTqmp6MGKtPL6XpFAcvqHEna5OlFhYvqj9wPstKSu
4qo5QH6k6Sk62zZcixBmSELQI+fRd1KFPD/LH6SpB7Emfnsd4PSbSg9PRko66mscNtRgkSIpjXSC
KSrtKIQeP/1hlEBQMLyxkuQB0MNjuiE8pHffiUmePo8uYFocqbupBJFirXx+D8HpZOFvXqiCp4PT
1hEsEvo4PUzx2iEO0xGfHl1RaZifRkg92Uxa5ftRAAoqFs9kfoz08an2y8iN2HVHKzyqjXen9W+j
dTViZbMDPiFmFJA9tINjp+CAf7W8M9TSvRJsP7Wzi2EA3fU2L8ZIphzjBaNvLTWTYKXPy2sp9tX/
21yQfKowzIKjRMrr1HxuBe8KAYWwOON0QFyekKyeRa2s3yCkRM6H7LBebKcZV9NHNBvGbV75GTkM
jZhKZYZ8V9VcjqrO43T/CqOKU3oc5fjDKU2YSWdNkR5FxIqGErjq9h9F0JUHNNML7i9HlbNiOf63
5WUbTyS91b3/FRl9rUzEvEn8HL55x3SXrQgf/ag3SC0i55KNm42ta32sFrUOcULq+ustoMzKK2qM
xZp2NdKhqXLz93WectSOXAkEfPmo7oqJyPtJSRPL/QsFLq6MVIhjClSAM5NrENxymoUuNZcokhLX
DqtP/DIpIrY19MufYJQz1lNmAjriCTBOiMIDUQqkjTLuuB1cI/X9wog5hWhdMOA/Omc66fcF5S9b
8WOEkHmKC6uHm1JYzXO6xZ3o0qctBCCeoA1xFUREtaanuntRxSf3g0dbXIGk4wJrlQ/PRMbVbyG/
ox2fu1yvyHdMrPHqyuM0drx74JAA7hT5cxM6DGooCAvESQXCom74CDDbribXVW6uL2TvO/2Jn9Sg
ln7ndfRouOjbFG7WcV72Bt6JORuDo1COKjX5wm5gNZUVs6bakU9tQaXeShVMoqkOO9VdH5Xnlyzi
aQoaj7PjyNbGcO3Jn+Mvl6mqiT0U5FrRpXH8SJqAQ3IBsv/HFH0qV6Y/rup97KTHNY5343V3Q1uT
SmuWHayXG9cKtEgGFxined8nCfZuYl/zySG7Q07mQX9gR79gIlg3qLoTxQ4oU2W72b/Xbqvph9IM
P/Bkb1CDxk7+7ZfBqBoAHDzE2Oi7BSNzBIRTRM6VBRCIShYRyfqCBKxKQl0J4t1REnvQdp4fBXoS
mXC7yDRt0CMN8f/98VMBm82vqTKt4c4CXdF/8jqK53UHWWjC4GLHqb8l/1Buo5bfmcblPmAZBDfb
k5bI9pqJZNPyHntHfqwJB9Nyh1u4VvcZRupMWaK8/X7EO+u46IUkdoqRtfnnGvOwgNPugtXEI/zx
AxKT0fL5708weLciDGXdlU3uXoCIHaG8TIF8FqdzBC7EkWqjI8/nHOdSYibbCNkPzdoXWMMLmvyy
TkvG6DA2jBagxc9IDHcrcMbcVtyQU29TgVR7z7B7hFUgZ4MFo2cwYv6d63+ZYERIV6+6zbMJH168
46qTfcDVH2bUEngqCCpHNAEyOVcTB4Vm+QdpzBVaDyUQz0mOgLdQK1CQXYkV/d2aPnBAzkybJEp/
Hu0hgTAzD7hI+Qb+4+1wXqNNQPpi3y9FuU6ZSdfxdmQ282L4d2Lyxzz6PE5xLcCwgiJsUs9N9dQz
oSIScfiPPm50G69LUXZ5s/KPBfEbDCoJMQtD9DYs/2kTi3HZi5QLcBvpcbhSbidGAFZa1AWV+0yj
wfe2EwD0Yct5WxF3lhhlu6CFf0ESNPHNWJYpXTqGzMUWa1PJuV1XwBu9ADEuBA5CaPrHErOR+OsS
u6UzVJeKizAmSWb3sqAwjEt3GEB/mP9Id+n3EqhhlwRs4lO/xC2WdzmgSGXBBdsDAPm+bxmlhlMQ
ZfE1yG0PPIW9GHfAxO1ZTotMFc3sOWL4o9/tUH1AgFVu/SeYU2pVxUluk0kJRSvTkOyNo2IMwjdT
0KUe87EvD0vee6bOQ8qqNFu+cv2bETOyGQw1mucuwv5pU+N5sGrnHOPSQ4H1OpaCXAliJiIGk/Bk
ds3pRFtmrQiLTrVeFtpwsWjyXq6akvSIl2lqneQXhef6+c45KaUnxZLUJ4Y3NVHgJ2NNk49kvYz1
mK0tJXEmTfmMEbqqNbCNYvFLTkmH9bCfmOENbM2Vwa19pVBD0xLxg0PEIXvVTqB6Goo8WPppXTgY
Lw8TSvscc705vGWOOGVxwhuQtRqJCsBE85a6rcCI04A+OJE9NzxkGopNqu9Bt/m4K98LFrgbuISm
PY10CWa4sSXgPd+8d1HjAWSDo/4kUdTRL5GK1SQHl0Mgpkc3R1oxwnECZKj2kGZAMuJLJ9t3nud+
15X9dHuQDLX9QWvAcTS5YbYD7AO7JSy+buZ90JrpXuC9pZl/8RRbrYiW3aSuyMd5YdWY0u45ahtO
12SuyvzPOxeBeQukGbOFPFORv582O8DQ8aTL8ERQYnoBtM1LPYwbKf5ThqtURFVs4ALeBE22yVMA
aYhM4411+hD298Thb65jIr20hCVLLgk6N6GFz0MZnb9VBJmI6vWMfcisltMebQX8FT4U9FygsA1n
5+K1M8CzH1lXov1pYbGFfEg1N+KHS/PL89oPQYsboUSUFkd1VQD/63DkL9NOW0h2toTNmyxBzlXv
ziKy6RSG1gkyJPTIOM/YuUGnSUnzvJATsNQKI0zHNB8rpSCTHPapCohJC0MHgmv3wIyKMqzofLlT
83VRBx85d0fDDedfVIxsJ4UAsoSedBr8XNPNg2bvvFDKjEiqhi5zZ4wqVFC34CewKziLfCpKvNcG
xIcraqn2vMWqFnH62zy4yQHeERMbeIMuwft0KOb8soICxqAnPPnH0f/EUFRbEKtd86BxX0UtMoug
HsvNESwimiB1Es/rIkVbNm4UGyxLwQwtV0S4YICvtBISKpejPTKd/ONcOIJIe2K7HsrUP9Z2yq1g
c1e22PxBJkdq9Rgbbn9hpNvWP1fLVNWQ//c+UiqcR2Skiqh2XQ3vpRhUGlNtuqDzFbMOaJXMJetu
tdzaCIC7z7t4t08Qxqn16uvANM7ZkoIHaoOwuDVkqv17xaO75LoIIbeCO+D0wnjx5RSYixzgV5ig
LI0bd3Wt3WuuRK7J4lsq3rlmPSxi5R2Vcr5usq7wRpEGYlzz5tzrBzj6I8ePqUtl9dXrPlsdzT6R
Sop6bFK8it21lS1DEGXLCPG2wMN0jyE0ZwdlElbSgtEwDjQFzdJO3qqnZHaBO23AiKOqHg+tL3xz
pfT+7E3PvjVLIKEuEPpLbhS0ZXPP9KD2p/SGEj02hOpFpALH5sNWRj5+NY85CM/2wBHqciwGzI8m
kk3w/+hovsofrwIWaRsntjfEXnXgh2w0APFcTkTFwzTkqezJE5S/h4NDc85+Tg7TcxFQOtbV2wwj
6bhESUv+/plGBND/4EDMMp+9TgZ4u+Cu4M7Xx4Fo5vqzE0dCMD7ta9kGMPuIWWoK8OAnBZIMbrII
LTCGbcBJsdNDGp3NT7s4hF9uqKseppufLVGjzX27kQZq49bw6cKHvmXtXVh7B6NHUP/EF0+825Dm
p5B+MkRtXsdEc3//D0VWC7ESEstj0VMfy4ZwhgA2rPYk0lWMyYgRptIV29d+d92B8UQZrOQs3+V4
0K6nW/VoDmRa5Ck4mpYv8KgkywngxJeyOr62S1ew40CN3v6Fx5A7nAuWcELaijKuxeQfv+71vTII
muX+xPbpyCnUac14noCfx6r8STznM8qNSrEAMaJ+3rBQMeFeEqPkxE2BQ0Ev91pvwtTLw0wgGWWJ
Om5B/k7uEtsOcLFAq+77ci7FZdgb19iqJAPOvyriwn3oI3euOR3AeMa010O75m1HPLYLkMHHGZIX
rP8Uj+MKnQoQWKDbo4gmfrq9UDHqNtBfm5mencIO7lefl4HbZddC0C/+/9lvJl/Uvlft0AzZgvim
aSu7C0VEc+uv4/lUVKyNt6cJSI5XHq5VOTDSFk3uvJ3gn+EXebfEgEobsXVnlUQOUdmCokQ2h1Kb
9J4s+H6jNuLWgXbLGByAx1IjT0SNMtW3n/7V9tjJ/mNeoj1udPZOXnS+Meo69k72zy4gVoKvCT6o
UQOT1upI/7jChTHBbvUhBmaGoksBqPYR8GjbUto4ILJiVFLj6wi5YSJ6jB3mguO2nwQd1ScwOTcr
9pYT4wrhcbjS/Rj5pZkG30jV0x5QALx/RRsB8VwYyxHI+H8bpOfaS4PGI5U9g/pDi6qTA90Fpc4P
2+rJI+UrT25Fh/Pl5xzhCMetLAzMGO8mlmYwCYXlLiQwIimxHbHxxqGnlcxYLm1LF4TRI7y+Wsj1
WNUUWYFGnSufbjTQ0d44lKs/hMYGsZNXuxllq5CKoNaW2Yfq+XCeaLKPPWPghNmguD7Zq5cnNQdE
b0xbGR3ZbYNtKJZJhTgPed5gnYozmYJt6lWCtvjZ4TM/PEEUpd2QNhMaGeNlZsmcIjBuqC4FgLfA
3BrrwTpSoKC+Ws7ZiV+nAHvSgjBwxanuIU/v/z8gk9WfxrOBqVlFSltopri4PyTxubQxe70MmluN
p3fVoIWRSGrHtHNp+HFjOqoTNh1z5Mwc32XLGqZnY8KpC0hIVHaYVx8WkRZ2t+e6/sAWkzZs7HHj
hhlf+LATCOzcwyg7dHiPZi7nOdwxgAUWuXnQ66rVt0VsIlnP8R7CTmAM6LppnLsXtHygjPO9e2LU
2LvA+J3WhKoybWD2neHC4Rlx0gfCYHSkP6409snsPkbgZsO9mrT9REjEJaQ1X0sEVoWUlHZhX+7N
6kgDUS8Lw9oq6tFJm5Odzj4If3X/9W/aqbKYqM7uYmUYgBhCil0H2hYVjaJ5HztTjS7Qkf0SqMAN
4iaWyVv29QcEsSZOQkyIfTZ9OKStPFIUBKqyKa8DVeC2TEPQhfekIvChJXZ/Wn/3MfA1NYwR+k3z
VrJhdpbu1v6gC8VFS6NjuP0f/83DY4XBLJ2k2xoJIwM/v3LvPoCl85jc2Mig12XmJWfO0PbU/Be6
RjjGfOowZvIef4EYosa+hOCXEio+MJKShr1YLSTyvfdmCWcObYV28wdPHFpJlbKExT2aG59s0GEF
2k2g01a5c0z1d7LcOk66ZO66M5AF7ylvPzyuUlCw8cz+9KPv8yHOTgM6t4F5WM6oIFVq65nWquSG
0ju+YvGcdmOYlDoi5yNZNbLlXz+xRgqIAbXc/MIvRfPdCRY9bBgx6DWtI1rnYlZ59kzDrOXJvzKk
UNIJZjGkjbFx6xb3X6eBFRmJpiRx53laZr85BPIvaSXsUTdX9tctA8XZgdRtuoCTLU0FvRWWTZel
fDNVdDbXgcKy/ZMEk5zxVPVb0HB9ipcxUMARSem6brwgf5Zxqgq+Bg7h3V73G8S81bsteZXksQZL
TxS/w/cchhelZMnhiUIfwV/9bzzSfQK10/nozfI2U/Br+a35I4CnXKSuma+1Na+n2LtdhFnR+Ivr
nKopHtmUN0HkwRl5nP1GvAR3g5CNasmgcoVJVczds9DNEIo67ANlQs02aqva9auCfT9ojOg/ii/+
hohJeGWmqxozPFz8Z7E7B7URzOFzoOyVMMFXjXRA9D6aP0NWcHA3DjSXZ5kNq8i2uSnUAGpoDsxI
uG3eDOS9hXKeYegg9phPQlsgWoDlTHYeuq8Igh5s7NLSUrUDTu8smAK8gbqpgfj3MrtFxvPRLSuz
Vg8citFZ8J+MLMCFsvuiz77N+H5Kaes3qgY/qsJPOhVHapLgbnrjmc6+2ZpvIsQc4XVWMaZ0lI9M
qd3KMqoozW6B8zVTDnaQd7kJcbD/bGSTubsoA2iCorXSgDuJ8Bx6pmWXHPik+iWDaTagHIrAU8hg
tFtkYlVfH+O5e21RwcgNsxRDHfzPWKlMITyZ2sDtiS02AIiSs6SveIqUFVxx1Qx5mvYp4+qgy36o
PcRr9wvvEoD+E7AhWuqpf3bek6BJmWJI7m/ep4QMaXtnGKF6dcNwbMrkmWB3WKCYx4hZe+DIpD0H
8Ty4M/i9Ud9N62voSx0XmqXWUPAIoWlRU1j2MRsVnMqTV1OlVhSomGTpcgjfqzmNn5dRlQCnLf1Q
bzPO7jZnadCb1VGYIC8X21+LucrbPvDlThm4kP/z1o4EzlZgK7zkMzrEu/hmG+0hVmF/9OriaXge
mJc6JefEvwbZa1HxmcwuNJmy6V8TBdXgpRtxqsEHciL3IaPeHzc5dZX3M6dktmXUeMpaTxP5t0nI
/x57kU9Ur3cyhQXd2ge6kygkx9N7Ww2Afz3jvIFzxNM1oBn/+6E4+cbkUSs2/ffxahUArDdXn4/8
T0Fh3cR70IaBXvpmkvyEK6B+8TuXblR0Y88i07+5NXkK5z1pOVM9+otNAHNWLSKsIjNys7W8s4QC
Rt59MRth3yboBX878Pu/JZUWcN8dzE6BwEou6HV2/zQla/3EsSWWZLKLM5MzIR7iX1L4YPWENeVF
u++X0/FmLGtVzyF5mqpG17Gqn+TbpDq8MeORraI0V4w2ImZdmGm4v3olpEuiiPkfY/b20ZsGo7vr
rrp/vyGt7sL1xJoT8BIyv8fE8JLiOxN7msoN20iB04+lNouuEmtyPEfVQjGoZHSEPUGM6iQrLZum
I5SQJSJXrD7Qxc7/eebNiPlAaxyz99drUXRa3tQ3P+Sg1OsALgqSBGmeSKof78f9HA9a+Tz2PVJm
ZjO+AVmT/YdyRi7eT+QBAaM27q1NYOqcwv1iKVV2nlXDBYQtKT0jns7YgXr+s4yut6jRt4WztH6u
U8JcG4AR9v2CO+AV04jxVngMxJoQjidpyELhK8RiClzlEIzUbGlKLTNd8j0i1RIkORwE13rCpiQy
1Z9Z7b7MYEFdShEmBpXUqrG9u+p2eKfvAEmJCJTuTB0xxDZ1dpGe/C58BU828lb0BVY9RcN0I/10
k4Zc9fEAO0ahI31WBgoCuIzpX1+sHntn2qx4XevBptz8pY3wOROnNMyinSHH2WRZRfUr/VtcKhSt
0tQKJdg05VvU3FIdPLMr8AfnqP1sVi4Lk9CV/AHMi6jRGNwxUyIS2FRtloqskVy+GWsGlFFGpzoU
2ZRpbxBhn1W6I87Xs5SMpj9ce7d9xNaIjBKICA7yi40iBEGniqL48sBx7qGnxlFzWhbbkwQNLGhi
x+aXFdwrpUOSyZwHTyBFS2+UCIIk3fzsHSzB0rdXKK1sfPMha7PZzCje4cGxA6627y0obj/UHVwI
D2Rn4TdKKMKjYkpbn8IHLz30z1lCzOJgaNUtmDsRvv/QYUosbpbrnnxWGJ++YJIzwUa/zuvndZPk
72L2miAocBb7wYFYi8S0CL8UFQPRDQR+MinVihf0xhBMqWfWwmAPniLFKEtmyfZp8NpguIUU2Dzq
K653iUqgfXMEXG/1H01SiH4UOCW4xwDCK0EWwBplvkoEQmKP+as3XEiFFDFk31hGREsZKfHf/OW9
hZ9v1Qds53kQqCGk/Unp1tD1GgA+p2NnA9RL3KMP1wRIe2jgfx5a7uUicr8CicqHoOopaWHcrMF5
N2ZV6XQBMGNz8XRnbx9WMctxe4A35uy+SMwsu7ll78TEFWwCZcaDiO8QVC47sAtKLdjphnu36U4M
Giywz9IISRtUFmhbYmYlSxlFuecV/xv1uiu4Gof0q+zGpKgROCoCrEM0SZ90MubiIwOLL5KhmScC
VuCmKDFEJU3SAypMe8IrQ7qukYevXBeOlpZqKq4os+QLrdF5l1K2hH0m2sCA/xNkski3lvut/8TN
zVkQrAc4wzJX90qT95igNGtODIrMRXSi+uUh9XPqJFkTt6tlT22kBlb9MZRVCAwXrzZhvd3dgVNF
WBprg1fqiWepRz/mVOLJ0saN1Ulj9zy0yJsSC5OclJlf9VDzNTGE/PJIkIikLC28NTZ6Hf0t2Q5w
pRDbSE+JLuJu4jhGwM/2Tq89CWfLEpu5qiakdu+rNimwnvKVQPhl0Dt7mlDcbDtOpMKxIuQVH6ba
Mh7aGq4DUcIyyPEHezzLQCSxhmjQEcyqEPNhjccFCj4A7lP115uZpG9VDETcwlHqYK0zz/YgdI6/
+EC4Fb9nzJfFEEGtgEvvQPYMjhF20NoV4J7zIXSFkW+fLduqmP5iECIVEBRHo6XBCciFVTKFT6zG
ypsOsmaWp0ZikG3xWHKz0NINu9WphVEVSqFhPaHxVVhE9L2qERiMS4Ab4j9c9LWQKV3KOtLwo+q9
TGxREXuHHqvs0TYcfymt5rbSQHLoslJBT4pgU6zZdZEM9LAfMMld/kjhH6VP5NG0Km2R/NvZK0aZ
Uz+gfRRAE3Y4UxFbcCnpQ2XVtoMNjYUYY7aAB8xk1+CwlE8HYuiSlukLq5gi+1PuCYOwz/WhGQ0B
rK2h5LCLtPK1lw/ZUm4YqYVX+yiAe/+aekEJfuUFic5qsppMLjwYizoAgrTWlt/FxXwgQD0nwXAg
zywSddNGC6O1aX7AEBIQg+iqzARueDSxxLSgvGdK/DNdKAuhwuDSniSnl6jb7CVzfyG5hPlFX/DL
UxS+/YkBKA7I7doscj7SEgkylkKwsHVs2+8Blth5w+eoBASyl9EXfCxnLQoPJ1BFT+DBen4TAnbR
Bjv8JLN3MicIT8rG2D8XmbBAA59zNApc5CazG8xDVJ6wCOUezgY+UnWYVAt9/deAnOsuF4WscnXf
f2ccbKTKvZsrYSj5qbRKLT+XxI5AxocxTM+l7JVedIi5SkViyGbcZaedvGpXlsyvQ77NBig83LDU
jlzv/PY5jWOOOuB659lqvPMiFG+u+x8cM+QNMrWVJrYQCUMrP8k5jUnOjE99SCIGHpiTHt9PwH1p
GWyshSpEywqB9T9XsyV7Vg1lwrhsHKo5Z4TiRqHdUrNBB1/bbdI2LcDwwRzumwYZQdJcdv3Lf/A5
ouqNKp78KmGEasyBAsB1Hp+58+JPwmrJAzgQCw/Z5A378AqXNIuOlzUfD3P89DaoICo9usn2779T
a7Y7CAf8XNPrv2n+UNZ7OGTDcmCNXySxDrFVksAOVSr3l7yGQnzEdou4pN2UXse0UVCTSFnczYfJ
WtCJetUY8W7qesahhUxk4WqVrEC5P98AfaT4FpbEETP4Bzlv75AECO5qmbi+Fbg1Pv6dUL/rsXkT
mtzblSqT28hJK2ixRpPtSNg1+KHG9AhqLJ82ZHjYkT+rXpkp6eKWTxIeLL/pMV4ajLk+a07AiQQH
W5g0/q4Lp7FVH3CDNSWtSLiO1t2JD0uyzuqrAxs9bShJuLqed1MKxcozX8UbI0OqyoDweTnfXJiY
MUZtG6dUx3L5sMkcBrhdLIX3NF52AJTlqwD2bPTK3wogKqAxY6TwX/oDh1qtLuodesClyzGadPUu
pu2bQS8qJdcOr+w+QyOroAuPfseRpVeftOs5hAsAaQIoXc7yN5Aq8U27ibVdps5gHZAAR2nDIf+F
JVwM08AR7ZzE5YZISFY/0KM8pdbdsyVCKNNBJFTi+2nD3flfm1aKmGi5fd91ASyR3a5i1F6soH/s
0yw0/iuyqARLOEv6+HEfmlHH37aauzP1wubyYmRAH8HhBkmSnFtAMAvJRx8yq1EKT6POpvYQuw0+
xJZaMBmxcVMu/4ae7HLg1/mGvY1rXrBPAnfDRVHNYh1li7scQ++NK9r9ocw4sXvwHE4/qy5CDIna
QseAhTIObFNNF5uBfLXxuDaQPBQ6kUx4DgOt77QRAQ54/SPLcAgCq0xt4IoL4THFBXNTxHpWsrG6
6BaDVd6GomWeICblM1GPkuTQHfKnBRAVnASLYEdrd13q1cXOXDvfOq5MhoMTLEg6IlkEGTmvOdKj
Uw8csQuFMGTS+yehwUQ/irbcKERoyoptYvIdPXKwbmymTX1Am9eFtIf/+u7eAJA1lP2SBmQ/UMn8
x9UaIHRmJgSO82rICrkqjz+M+vEW+SyIBietXlhPjVV3f8qCI5DkTpn+IVAJxk+mffHn0z0Uh0u1
AYpI4hcA0AWMn7UiTG/UDGPfa0gfjeWnUHlGgfbR2k1pGzvdi/7QirbZaN5sjxx5vn+lLWCUCHSt
drPbwuuCK+jR7tFtKNgjPse/coCb2YBDHiUfKiTFrC6vEUigxr64+nsGh6ke1LksP9j2R/gDv+bN
0fCtejFiKdSH6NqKJQWn/6tYiLxzh9J+Wp/Y3cUhKKDXKmYIZSm5ngQGoeTxStI7XM02eoKjYImD
Het9voYzYn3ssQV9ZquDNiu3nidtknL8sRGB+XsOSeo9LJDn9IcEXz8MxIcfcLgO8kNAdXLT9V7t
NxT6FBcehJZOkmPEFItYQypKC9V1AlLovkuM+yd8PzYBMfjKaOIzq2sn8N6BB6odLwh9tdGtEjKk
FJu6gmemTblCIQm28J/dNvM9OxupgVRoSrSTsjnWeftrby/fNR8IVxypLSz+QFKwxkurfqo5P6EQ
3pYI5kAbQ7c2gl2bx6iZvezfyXXLbpalFZ5jikWRZhBponHPVy6KMFIShBlJh3obLzxGgREv6FfG
8SKQEL35tpxcvsVfzYA/opQElC9M8RchCDbZp5rtsOPRWt5x40IT8At9kUHfXIWkYO/SOMmVdDI/
+cyy/VRCnX0+t85kRcJA836vkAyszpLo2Q46N5j9+rRW3HMV0UZoH8qt0MWoENg5cjgS+WF7keMo
W/+mlwGhmCs1pnhRF72wD52X4K4Rln2v2pvgXD5qlfusngC8wLXmILCcMV/Af2SqI2uIGvC1NsN2
bStZX7sUClXyqZCP6OpFSjSkoTKfI3aSP9D1co4by1yiNoO0lyLSBQ8w3dv63gUjH6UldntYf8r9
ThfRX1Psqqd0kOocC2ldeqwk9IMzXiVsOG2KtuWCclygPOxwhlyVUbd6f8JtY/lgjBZIZIft9zcA
Bnbm/u/aD31lBmQfuo4K9daNbuSsLWg1Niw/5G7ryg6QqQBKgkhNv3FxcuzHq4sWmYRCJFS2rt54
7Ulq2/CloMa3/yFw+p0UtSA3hYM9rCDv13iGqQA/MaPaEXtaEL5tIIzbm3TIG1hMCWyVhdGEpnyq
kvdDBTF/Jug9LVMg0ZWetnRvs/UzR1Xjkin+c+tWJHVR0BkGJkrJ86CRk9h13mADn6jV5/Jk/adX
8FUFf/b2s1BkuoceUgPaorlAiMSfrsUxJz7+Z5T0OH8VXpsi3FYxBcmHxEWCRHhRQ6ORFJuIiPmp
aNEQ6YUKFRFwS86+zgMOeW5u4gNpPlDGjamV8DaleeQfvf11wK+ftP06wW9CrjRe4qzJO0iB4QmK
fHwnSdJUmEqcS5JIkeZxkoEdO6gnRD5Ngq/JO2kpz76/x5Aj4n6qRhtpa/ej/4uQxRk+B2Tir+Ct
K2RpJmuknQRmwoMTnzbZ/pnxCsuJdBjC/bWKKDAeHv4P7SE53Hsjbw/Ot8EX4V1xxV6f2eegQ88r
liMEkEG15cq+w9TDUNvLI53X6m8y0ROCZIoHQtFkuuIlkOAG8vDygQkqRQaDaKD7AQvYRNKqerWa
oWkwMzam8nOJoVulzjJs/5MMRF2pj9+B08y+zYk+927ZnZgkcslrY6MXjqYWN3t7Z3GiZ8gEMxKq
RefFigrq0luS8GsnqaxKZNwat/Sn6//KJL3TtjvOBecA9j3HJr4ifPdS0DBI2ePwC+nYfG6XTJ9L
Sr6y5UXzicQFaBCBoncZ/pu/nHQgf2G05Qe7RD/eA1x4k+Nr+DdmhxLfs06e5MdTHFvKqQz8u9v/
9RtPNJPGWR9PNr3GI1USiNpbfh2RSW/gWZUhuLrtl6JSFvpg+7dVAze3UYag4bsCWEdu9nST+exF
ofOJSOl/91/Oj7leviOJwZk+KtkKwLXPWDAbarWxOzykkLZgqGat+KQf6to4C+X7x5CocGK3dXe4
Bh1JQfzprpvBcEyDU2deeNokJy6moFNWkPhsyIA8bwhnVpzXaxFJRjQe0Vs3Ou57eoRNj4Une32x
aqTX7PJh3axHscvfp6bPoqG2+mzTqUTM+cbxAEekR/oeEyqTqca576XSurLWUGEfNU++sCtL6EDL
NdhfLyoMNjGq7iEMcG/jVe7wDJQaofOqZhBYGM3NXR+hYdqHPooPyRIVApHFMOHi7J2mX9ivI+Sg
RKSbiA6bYftU4O/+xt3+Gl1Zs/3isQH63dPNk8/7dH4n+wwBCy0qSobGt4WU47fiNBQCkstNg+aD
3T+Xb0UwxeXA5HN0sFkPC7BOhDbCJhdpBeFMun46dlB/8LdinhlPFCLVumYaleh1z60Y10uPJ33H
BqYNJnyUIkCiS/cyJHiuwcq7d39ytmFysZV4D0bUwnAIjvUzT+4UAYGnLhuJm26O6vOYTq+EGH6b
gnIQMGaXrOQjDl5ulJujRd+Wwh4GRXBt7MUeOE1neD8ijOuJ+PDK4SVQPRHeWFPY9p6ipzsNlY5h
GUI3ejG5V0Y17CtAw6FwWF2AYtn6OJ6M7DaoQ14bWo99W7pPYCFIPNh7KqlFMcLcuC1AYvd9bIwW
LPSUk4zuoB0jo0Oiiqb1BLzbxwfnP6DkvImPWcWtBTrvDBx2JBMAfBcUsix+7ezLp4jsssTtAJCb
PYEIvNG+V0KIsisBz6U96ZqL+nq+u5DPvTUAiAAokd99DcN4mgPfPMptBvM+mK0ka+5fF7BMRMBk
vvq3K7TZkBJbeHC27b2nervBRC0MeFUSkjRe1e7VseJj+widejyyaR1eb8H9NGzAyG31oRNJok9m
UdOrXm4dJslqxLbIy5A5PLMmfbfcjHph0SKnNEU09rN3fKIpLUTipVEpvsPn05VXxmXyME1T3590
Z9j6s6j+083SPRY2n0qEN/8+XStOVLVn4TV+ZucQ2gh01narvkIgh+9Wzj4DATeN4aJNvbLEo7g9
yg/vvxdvnLHxfkkE1+QVLhck0jFpKjVcMAokn5fiFHc8gg3eN92yyrNKj5F9E/wvSxZdRSzpQ0n+
sKlH4WLVck/4nQ8gtnt1k1ITKvIEsvom+GsDsgTnWzsBUjpv3xwRs0uvIHqQZx68dkFch0NV98fG
I6h+aIklxZG8vEggbJEW/wWdSV+3rLuneYPquPmjVGb2BNOApZJjaVlSX12sK80KC+6KO43yvzoj
yz52imc0gCormYmU1Mrrj/Q8Ebehy5iipWNuPp8u3auJhhX73fNreYK778NUtZ+CnqBms5gpM7hU
Yb3s1hdNINgqH/bDnZz3N0AFClNlg9kF0m22qurQ9vQYx+PZO0OEFQpG2n5hzEiGdWD7Kln9Eux1
FcTgiURG5nLw88ziBDnTYsdneMusvlezvZAwBCmqNh2QVrKe3b9E9CWM8Mg3bda5Hlf8dYzgdEYK
iHd8B9G7Vf70De1firjoAK8UBJDtmAsh09HoaY349vo2zQMKuaRcwzTigVkYA2nUkDww83Ny8Us1
Mpru77Ydr1eFU/s//qe5nQz1qEw2OVy74i6rfl3m659gN6LUMI3iwF/WXNIUs/7QbKgcnV73cRv2
pKXqwnGISxQL+qNyNy/recaEnmTkQbXiRIey/OdcnSx8Mo/9817MVpnIuBxl5h2pSGuF7LNbe5dX
ZmrDxV9uqDxf2tSfU225WmtPyneVUzQyPj+sj09Dqu6bm94v3jgoV/IjsuRXdXLkpws7OncUsGOE
65s4AP+Pj8ZgCTD+8pqJpMz2BfuLz1EykhHSokODwYVl3oQyHrnu7C54wLG16iBUSqgA0Cu4ycrh
udZJw0h/l3IlF2ULyp2MzptyOoKqTh+9zHyRYBjBpinaeV8ZrXAcV9thuspv4I91Mr+aKil/eQqn
HCkuucQdfqRsseGe4heAe4BEGS8LE2gblOUVjOfDSMFZ2py7hWDzJuWto+Im/foW1KYsvnnW9Fpk
dAApOe2pVOSLhrsutGCf+R67tx2yy4E2KWni0hDGj4X2peuIl6Y2a/S2YEzEe4Fq/kR8RMNih2SS
lOdFplHrIx92ZvFA1hIVgBCGgxuJg3JefOwyk/0qELr87OimaCr6cidVADU2hGKqPiO4/qa+p7Y6
0A096nTYQmRqrlLLXiWeDgApUjHqnchG2t0RWbl3VwFqgSsaV5IFm5B4esKTIEVmgw2LenNgit0+
4QbZJUEP3q2fb5O4PoGNs2sg4/wA30K6riBMKSq8G31xkkQ1L9X9LAlRg+4qJSoPM05jv0lBGRur
EdYOLm0NALRT2i+TAxWyx+qzqJMVgTmPVTIDcRSCLLE9cu/qMOT1v2jssy6uN8vGPWgC2mO2X+8W
wezOozdpdojTBw5cYhMVD9obQgf8SX+8w524qO1CqmQG8Rl5p6JnTEo4e5EchYTIRuRb6OaKNTKF
CUd98knG0mRvpSbDROMHtXIPcLtEiMOmy3+1v4q3e3Ou4DgL9/iGwuBd3Fo6vkjfCrIQqZ7F9bYT
QDO1z41vGHgmxqP89/OX2vzGo0EoKPNyWy7YY/Qs5+4fCYyFmkI3tkU2RVIcIct+JN61Fx2inqSs
vkFtWWeHYCAz62OxU0HE49zIQUS9mA5/1KBOxROjJEoRnOGGCNPQHnAggiwIMmGVIbND/Vv2jBVD
7zJJNaPg5NmnOI5qAJ9zEsV0WL1WKTR7iPHEg+2f12X4OwIL0DKPlNiA8zpRxdoVSF4xzLC8/jjC
256mSUDk9xyV5jEEGs2b9eP5E9s1TvWyn0z7RGDxYWr1UlHnGQowcqDE+r6lnqxj0idWhFleZl8C
Za+AKcqguPcS8glNR82itihVohY5wtdW6aYhghz9CkOh5BLBt+W0xiBXGSk7xZCCsD1myupoU4LE
SSVJmq18cw0DgcnDrQ8061qYrmdBi8LNtWzckOgxBGAOHpMJul77F0kAoOxkCLLWJeGDb/7Hbgtf
ld9cSb2hPC5xB2sduas5E1AaFY2h+ayMbxbRxQa0gCEh6Op+055RQINPS+kGM5c5/Wb3OIQp3vbH
u92GudI1fBUy+nmQ/OfLrEdC2qol/NMR1dakdFQBRY7Bw4l1NcCNOk8Rb06zYIWuRyNBCmXCXY6k
WeAWtFNtk7MLv5O1IAqOSU+SnMp7S/lgnhg5CGfRmcwCW2hk32ukFxM4UfBU1z2JHsP++lw4PhF2
C2wuVEG0MWAj59TjmYTO2+pEl79G7GJ6lk5HfzeKdIsGC6u9eNaLiLKWIVZfp/Z0i1e283BI1V9W
x1v77hZYYhJYp6gVXSg2brHyLuMpwc3hvG/lpLVTEMXoiWgJXJyQJpfeV5/N6K5bo5equ5vCGkJJ
7PGZAgT9Xsni5h3qeeCUdB7gKZLOPc4hiagEaG9UJiDn+V4WdLsFsSjnItI0La+uFT5x/oEqoKor
OKTCJjgLQWpC/ftzn5QxMJARNpTor1f4yPDgqQ0k0ddym5HFz3RbGuim0KXYUXoLBp5t+kf5ergc
bYmh1Bq+1by7sAsS4nlv8gQJd73UbESMHfW6YYzLmamIt41vyGXDIL1cnv8yQ61Q10uDrv0xnayE
PKpMaIsRBR0w+DVAFbzPlFtu2st5t3uxoKRdXPiIqmxleH47oYN1DMFim69ph13uz3PedhnT2+u7
wV3So40uNO4/K5p8VA1WhaTgvXx8VV5DXX2Fe2ep6kErujKtR9Eg6s+T6o9rElYF8RH2Xi2rSPf2
kWRsoH5bDziWIhp2NsO4qPPN43iv1asqE1DwA84ZV0XyJCX794UD6RpZKwvRTvW+atRbOaordxlF
grmEHQXH+IWnOOo0IIrdyAX6GDsi9T8/TT8i5t8WYhHN3NFx5xF5Qd7saSrjbnwI41KEG/ubQWdZ
+c8y8ywsRqJMRLMN2Zr1terQPASySsjKdT9jFS5VM5Ay7Xt6tkOWklBV5fXGPgHTl41mzXMuaD5i
2+spR6SRjtrGfKuA3XOuFHDtjVGXqJuMsq1dGoCrH0fpPExOvIJJUZRZTCxUKl+AUeFW2Sau3oON
wKhj4sO0LBhphPaj0S8BaIUaf77/XveVRKvTNVo0u/YSKEZ14i6LqI6b7I1pQDCmEoqnsfDCCHxp
5fZ2GDaQHGa7ltCAlQvFr1gn0NmwskZeZfcrqOwRTF47aEk6u080oLBSRZX7epVpPr3jXShxTHT/
Ohjfwu8foZb4EZOnYbeDY+/IrZM8dbGZv6r5wHEsmKI2WI1G4fwg9xa3f/jdFcWjPLVeOeoKWvA1
j5fAJSUFodJZHPXCD29B6b7yewFGAWlOerFQYu0ymNSOR22G4Xk1Fj21dOXQkN8qxdopaAQIjra2
LFbNi6BXZ0t2nKiYdM8dlRDiGz3PfpALY9JvSsCEkFvp/y75oAzMbJIVatAAOMchi082lgytg2nc
X7GhgD9TOhpQsmqmdqlin8f7SYKjsRhPhLJyjO1wOiHnXKWg3UhOmcGepIMnOfs0lV/eXab76RX4
iJzilat9/knxF+h3TaBzCnz9dgkdjQRHZgNloWByLz4OiyZZIVNy0SlFdk9+pLDD2hOv/KRbQLuv
yPJzqN5tGTJIkxojZhrF6AEQ/hDRTowwRbEGqcowmerr1dM89EDvEwD0Aq/Iq99vGifiUd+8jtU/
piMG19rGaQ4HXfh8Fr8rtFVasruiIeGmvKR5/cu80vvvLNAhH08NqvEOTSjdlSb2f6cvIUh9AYAU
fO5G9pgJ4QhdNWolDzW5Xo5S3cQQIMonmroePb4tq9RlR9arukq6QPwXaZWkcgg0X2QLHkreWBh3
pmxFRKcvySdCqxTALE+RbU7oGhIvwOOLSGyMu48aNwH9o0bArgZycFSbyKQ4YFbLI344dH/eKUqs
6nAtAC9xNPnyua2IzAVvXsYadZao1q7Q+7LfwVPr/HISmNV9xDFVhLOmNhaaKoqFl7hWImSNfX4n
18Vwpkr9sWW027euYq/pAFZ7OUppmVqmoF2HO/bF7p3ZQ5Ak+UXmmmwDXFYU5lSYDYWWL0AeU4vK
0eoazgjoku4pZEAmQs6Fz45plMgDTHAUIdIWo6cvUac0hmHDHHaUei+mOXKG7XlIeTkX1yyoSKi/
ttIL2DFctriush61ytmq/xXQKEWYN8gHHX4P+y66dvkfcLC7qpqott6MdxIk+v9GswWZqt9iNHYJ
/zArf9MrqtcB1JvaUTAv+bmU4fIiK+dx5iAONiBjbc75GZuapZAWgpCTBKkaXGocZGZHXJgh6gob
ko0I7sSEIu0zhZRmiNtLkwFvZ4NW71WNzueuWEZONSE6Hv/V8uXFMDCNU2CfCIibNGsW+2s0KikN
R9k4CRcjv2C3/LX/VRY9W0Bcq4s7/WQ4eonIDQzu+XPBD77E/YK3KP9n8s+I2Uu51LLMVm40HsFk
aS/ruLbEcODlFVFz/zzDxeJDWaK7T7vf9+MFAymeU49SdTe5Gd3Eby3TGuGc3Er6Oo1cXe3wCrcQ
Z60D9Fdlh+5oZScw1f5uaF5u9mpN13idlD/QSrxkF5HynvsJxw8AvBoUmdJLpBTXSN1xwDDGzyQf
ltbdRULiWkxdbMZamTViOIwBXpc1IzFrsFmCfU8fixfHJjS8WaFl0v8ILqgiRRnlNVpSPioaF3cp
Y7ygPIssGwzkSQDlq9V6Ld6dxayEUbfHUa8CFWOs53gFNT2SyzqoSpfL4LRMELO7VFdfdcBK12NT
s3edN8dela4H/EMoO91Rlknt/bEOZUn0t+6mMc9EoeDvB/aFvjgGN1CqOlUnQ2AGbuokrJ3vKh3d
jOJcgemDCf1vjBiG+6wDbhfrVyDVji9VfvccHmfiLVpcOUr4wuQlTdI5GM6D+T/AvrpVV1lW4ukf
JJWHinUU66cF+q5yzBCs/dnCGpioPugcW53WiDns0m/XJzRaAfooHH8GE753fCHk5+RXk5inoe5k
NqoI3oHTR7eR9sAz0lREZQtyaNolnIvn6xkFV+W7SdY+1bajecxJWXguZpxrjRFwCAe5Vqzk7wu5
2r6Zfau5d7yAeyjvrjGdMqAI8t8PFEZLT5yKx56Gc+bsOFpMJcGvMhpC7zXRh6j/PmP1ZnxRxkOX
COxyY5v43ZybvwLoWlH97YZOfhvv5OQ0xV51hG/pqdHb7WLnAEAoX7/5vtqx0GWujE/Dc6rr9DzI
IIAXYYzjXc97br3PG2cSuh8rc3nCIbbRD8mqgvI8dDuXuLZWS4AxX06KloOkitscE0u0BSmhzqxK
O2zmCHBj59/NGqgJoG6d5N8E7F7b6K49/L3AgXCQefs/cF7AkldfyiiKaa/0zSuwx8gWte8JfwiC
X7qFz7ioSt2Lafzl9UXhSje+dbhkdWoBLN8IvgeI2S5gxVt2jVRKz6QCOBrkRD6zjsHYzSEWFmah
2qfbibdzy5Tm2nSajwfgc//nrJAn6LSDW3Kt2/T8f3LlHB6wEbZWhjhBn00aZ2qp/Yya2rRu+pw5
RZegVGIN+LexKAT0m945nCgz+XIV7Bvt0vrGSKsggOdDKd6+aQK4zCkpszm3ge4b2x4H9Df8rYSA
M/7saGfnqphbESYEHiH7fcWzJyKyJd5M/mIebAkzc42UHPyB8BWLY0Mpm2JwY/yKLkOlVducStki
ggl00L8y9Ei8BMBmGj1tUfFzbF3yeIbIzUQGwgXqyoraDsFLyUocfYRrEEpZesv4JAcVEB0TsRxi
sd4k8+FwzC4lEy7OYr/JQBkVt8ltByKPPG3blulNR2/JrdFJ8CkKIZ874IPr3Ofk9tMB+EqIzr+D
NkqcLWOmA6fT4gkoZsaIsrbre0EGthrpftgspNFHq6YIKpJi69NLNHUb1ZwyDAhd+B7kDCK/5P0V
/upx/RbKQnjxfAlT8GX1KNeTBczBEMZOuT7tjX3kwJiEU9Zs4EqajRScewhTSTxrOxtqtw462yh5
Q+HIgxdWTjZPyO9lpgirhjCfAj6BOlRHCnhZE9Bnybu5D8TqCEKl9H7NmhpC5IXxubxq5uonAk6h
DKuspPPwdP3Tpr+HGoXUn9Ioj/W26SK/MldzIHbwj8RbO37L7rxFl4b4/yQLCyMdpWUvOaY/i3xE
m0+ICfYC0x2aoU20eYcfkynNco6GPnsQVxnHkzlmKZZnuAotLuk+J16P5Eg/66BG1UGrNjbIzEZC
wvMl2IFijnLfmvMvUXa0RK33L4pGqbBRLxFrUo/jWCrRM3ngi9Kt/5fGs0x5gIrK3OjoE5eemwp6
uV6x3Q8hO88JRtMl5oikrGLSzv9ncKwwYCKqS4Y1jKC3uSOH9xXIbvUGQJFHbHniyS+UPYGHJzA+
din1JX0p7K6dzVCfIJeFsFYByipRu5Vg9Wf8bomnAe+JJR+R9+6qC5smlHQw+j8voirUhl1p0Me8
Xh1/Un5hrfTDnG7pFNH5M20czFtjWa74Hxrk3NG3sH7XVQp7qNvByWABA9ToVTLG3MBBBBbhRMZR
rzlJRSGtOTB3GRnIhlIWrxi1ALeP58+uIBGw2vtG7v0Lh1LC5snYqFw1Pe0eUoVGKY0Q1wUKo5Rh
mWlxrdBW9LXKa/ZikQ36S0cpHxXnPOogTJ0fkzUFMqDFazQGunFazvawdfQqZqLu9iwhpiujQiTE
uEUWGn5lIhBunyNwheo2YVxGoiqez4KAjUdsE3CyIM+0zGSUbclC8CnM1rqchhV2D8TtA20am2UV
9AL++jaw4BRXw9u/xXxxZybnpYFTXUIY8ihn9WVXfuDQPPTlXYixORV6E7moT1/LtnksTBuNlcU5
JQiMz9Y2Ap6oQDJU3LiQ6gKsUujWgPhBtzHq6znEb0WBtDSAzGquW/npJ2ITaA8ZDgNnC7dJAe0u
2nQQG3bjvpaXi18PxjAsidDVVdRwDDGwfQnpQfCgTvoAyGtiVaLEdBk/vDH7S4nN5jXl9UjmTMW7
TKOr++DllO+PjDdirZET1nG8YsE+1vRWJgGB97X1kHq10iRNV7dt5oprdDYgN3H1n4lx8RoHsmvq
w6W2Y9GOaWdAFejKQETKmvE6NfbEhL0RMCBfvqEAXRTOH3a6NQ2fmWwVQ9IqCh6tibLNKTZ1gJoN
0hR8/N/WuoUX6GCEdkK5CWZ473AjXwg9yyCWH75sJwcdnWsrCl68TIJ7yvgMGrOj5Jos1Ia0l8We
UZj6GKSiFaYOg4DD9l+sc/4n9yAmz/xbDvbkSALi2/la+1HArxOb3QwEnezw7ZmBhVBBngGqkZPg
SV+oxsoo8UTCFAWtSfka/izR4OcdHtoZ3BrxU+RP07WSVRLJf88w1GJHa5AHBR3Dezlu94Ew6sQm
5u7hdI2jq9cfsbEIR/H9bXSwn1M4/2Omlscc4B8i1WGbul8YCI0kyVYvO2jWh3aURWpdC8uY/5sX
BgbZGuvVaPZt0pzv0qlB0LaebJra6WnD1iqF+Vl2krjIcBESIQgs95SKLIcTYI0Hwj/KYOni7Ulk
KfU+J0lUnG4t813WQJ88oDo+7x6tZm6qj2KYp4pkt7K9On4TGGCcf+Lrpwi1JDXh97Zz+1ZtZpFk
WW6+9yMZxww879GQb7HuQEUm6NVt0NSkJeMaPOhkzq5Jn/xP+x+0ICkf6ZCaT4OSPREdXqog93Zk
2Zf38n9hSalEaOKdGeEWGW3Irv1zEhIuDH7AqK6tl+xRqwRXKAxavrUkjtyKUXqcsvcYp5mVmyuG
HiA9z57QgjDkF5MvyJu4FdlKZazN7anRryGal8+OXsqG4/nyc1oUkN7arAUs3ii83h4WMM/J+8PV
dVMcSmuZWBE4M9jNFtFbZHzKjC0/iJ4ZCbZppkc5QUGiQPaAuKSTEBFh7O+L5FFSol3qdIVM19fD
nyF418XdIRS7M3Df6ta/deB5XrDxz1J5s5MiyblpvdUddUBSe0/HKTPbjtiyiY5Cw0ZLnQaxg4bw
NpGh63CPHDr8vYvUxuY/61748/cuj2pEIScFY6LlrFIkGJpY+Vgd5sRudcx04znagKNC8m4U8mVy
r9OhYW1+/XLH6zyiny79hGfQXJZKnewk17WGuP/ecGLJnTPJCNpR2bdbJ/y7b2YN7EEH7iClbK0Q
l4b/IrVUyXCpSvkWw4QdS15Ms1BHHBjPuwhaq7okscKe+Munyd/oWB+wdT6U88galhExfrOWq7d2
PzoM3aY59FO42fKf4NAhXBCE78B7RNOmLQEdNUX+LJa6DYVBjxviCiV/JlYDnxK1bETI3Ldw6kky
hbTuQ6aRHbg5C53m7jZBUjGrxYWa0CTvEi8RiuYewUbzTChh4cerHLzBuaRnIPWkSPgPyDcTBIa/
0zKSY4mEqSTZpROrR9G1Eo8BS2GU7eDL12fMJkmTtZOJ/xuaqgYVoIch3yOQ+7lzsn6x0APfozNp
3MdhoA/66a+KQ92fJObRvU2NVDIfPNvaMMvTTWpFKTYVfOvP5yb3vTJKpSc0jb2CpCTObo6bbh/7
tqNQIE7H5Q9l7MWplxtJeEmNnJIaJQKYU5Om3tRnb/B6jeSdCZWG+GEAV8JjK1WC1X5Jo1GUR2qv
yPbNbvB7ndJ8sQLD6d9/hL6ZZI13rb+ytGYnAYZSZr1ZWUpB8cs51huKZBmFXX7e0yjC8QTHrfYD
xR23PPHfU07pP6F5BW2h6D+ria5K1n3lKYNfEml/+naoT+Hn9wQbOvHuOcFNVF03VZydICzOhrDd
e6Nk69e284VWoyxHXY/ETCyvk3sO+Q3EvG/SSDPeeH+UgQ4AhWssTBj6+UjsweQ037DKBB5oIauQ
LR4s7ROwXbIJ7pxntOXFlcXd6iVzCx4hGETEZGekSZGcYQOqYx0fGQh4meJ6pQdUM3mp8UvQUsOF
k7d951qgwm9U8YRNj2eUiE/n4TXcbI/NukQB6pHoVJV4ALswoF0pkSY7JDWd0XjKVyPHGsKtHinv
GNGCPiq7Qlem5fyVJyOJpglwsTfs+45qbw3lchp3gysijgKXA9tEh74JyBEsxRjdPD+PuOZR71J7
ExD9p1gtkOPXFC2dtCpd2XqvfwZfADjHzP9//H/fvP4MxfftB/IGEStGFB2RPVjssix0KwLqdDLe
JQKGpxGi3iUQeQmpbI0x5HFqQ9f1dHiyesNrYlhWNwS51mwQ9EzqP40MMgV+dzc6YiwScm5w7jJP
tzbEzo6Tz6kuSE8Glu/N4nAzE83jQUiAh9eY/q7glDxagAM/dl4XYktYEMuv3D2JNwk9LmhKbISS
G6Jc3yQrLuuaH0RhXF/uT2E/Yh6we3vBCVovAkxWpXrlgh3vc4uuVzmUn+5bVqbLR4nhFgnD0jh0
ZkOckSX0jKGKoR6UWnr45DwudyuOXauHHPKL4dCzKqqYfmDsxLfjEm4bMT3S91jPM+SAVxG/HoLZ
pVaJTX5ATsnTWvrRXF+sGDlRDRKrCbE+QIzI5/lRR/+Y1k0Dz9NX5txuOlqzJtBidqk6lYo57Dfs
tfzqe6OX1eOVqv2tpu38opJ9Gxy7fQhEjsi1Heh6IPycGsHNwa6EUAsV7m/Hw2YFmgwK6y1x6pPf
TRLmotD5H8zLFUKExXN2hgycl0+sugHHJa8qfPDuIN4kN1D621DQ44/fwZ4Kk/wdw7KL9ZXdJdgF
pbdAaECOchVBPBKJq5RhkpgZ99mDQdC6Ecgh0S+u4qNXTPEe/c+zzIaxvmlThp9I/p3ozncrEp78
ktTK6oxNAgRYz7nvErgZLqV5HY3fLCwHK7IiF/P5YfHsPxU80oYesXSpXBNhNuLyb5I+pP/JXyK/
FqBsYBgx2sRxTA//d4SzCzxJ4seRsc7NL637sVU+UWTUpKMdiBtFqM6wamYno3IbOFsQeHfYxWCG
DdabbfMZyTfcm2mOmkV0erFAw4FJauIgXzAaa4YVoK1XMFUg3PC9D8bq+u9s2Iz5K+EQK3F+iJhg
hdXpy2uZXDHcwiG2gNgrwsPcXA2y4TXerM2NdUxzfVpuogaDrVb7PAGIKT44Bt6kdCjSnSrlEAkU
hpgtj6/plpQlh0lbW0kCPrjfLAqOtqea161fjHjgNm0E8/Tf7QAw68R1nziUG5QdgEVC7LUPJJ68
NJ8tsV5UpRV50HRmao9Vdi5atgt90aGeXwrI25vTpgVXFb1ts8QQ3bpIu8U3CNAOyjD9HuheVI5j
DugQt9wpzMPE6cB/zy5dU8OrxFcv3O2Oc1gRUipILazJNbxmVJbUOz7MElWcQTXCOhs9RFh8TqT2
FYPVF0ASBBaU/ZTmUQkFjxvE2lH6fS6G/BcUK1RaMRESnO4n7IuW7dFlU+WXxDQzB+hq6j4srajY
b6B7O1RHz/2geXOpBidTXcqb/EhLhjDFw3XZiB2jHxdlzNRsv9bUcwd+AaC1/tLfpv6WTXnvWEqe
JeBoAmetckQMqTSbW8j+OAv3TS0HXlQgosQPPEi54Jt1WWqHh13kHdmvKM+npMgbyKL95jm8rI9z
0URCUKM8w3rsbo6HUCyWZhR3QXN+ziXTXZR+q34v+3EL44WiHQ1pbH6rzNuak7aWo0f7xcS+RcW+
LpE01vra1/3MpgwXCREMa4fhtrSFYR/9T525pNXwTXNJXlQN7+nkszxp0xN8VnGZDlpSnF8hCHsZ
I5RrqsWI3wMe8+hC52HYVwlpZqWp1ehmyxEBg+ahHDMekN1Xm86fD4smUe3MIZuddwYeKAd37OsG
XufOLdlDriQ2I0t5UKQRf4aI6s6j3PPHOO+iCSuECrogLSJ0h6sxHkipRDsu7EPzLlKFRKIH38vF
lsJjq8Vzpy7Dlup7MmvM30DH4H+nPJxQ6phiO6U5rrpAppXyNVr1iOtBkb2/ZdBVhvxY9rnkB6tS
9mI0CMAtn9pJYO7DPT1JlopsCKpEfMAvcZ6D/nYRB8sfCY2n0h/6rM1l3nFJ6Pwms12hZ0VBFvaW
UhjQJripKaMD9PqqP+LeP5FfttUQMxXkrvKzFVt3hXSXaPuSQ2zkLrDRob5d/1kZ5O1l+8Ej/170
mzDwScFe1TAVbEgFdakAvgsMiNdP3N1ykCAu9ERLxf/9APyfVnptqn5/weiVuapTLNqdABGZV2O/
EGt6+xiiZYblcGhBThnweUuGuF0VhAhQJBBKhGd0DxYEKnG+Xh78pwHXgVoE+ATIluQZ6kpfNC/w
HGj5TcQiAt7a8rmxwnMQ8iGUHyNlf5x7IkwPAcwLB9LTFB25AnGPBbg9sTkvJEdBC+2KBpMRuUtB
bAmRrGALORygnLBRDGkWQjjsZyqJMh5o68tBXrgQeqSPz88g9h3m2QULand5XlGwJsC4Q4yBkE9y
eUiipZLFdnEgyaVA2Bjm871jnKJZOWEcgne7lzjTnKW1MMmKkXqMUIEpqGgoxf4vGZM75wakYJHv
Vioj/ethC23w3m+wbyjcp1NQkNM3Ry2Xq6Bn6RDN4K6XA/gjdDfyLRGSkImJLBAQ9gxo8W9CE94L
X9Cmt6jp9C24xcHOMRSAKBzZidkxff1j9R3dUbPF/TpOytAGOTt3Eqs7P+5tBPMp6fv0SOpIsDuW
UFX0EYehglTpklNq0SwXiy5WfI0/VhScInSQxech8c7J04fkvZQzOTQTy7ygJJayqimtKVVX1RXQ
2b2lSR7GQ460aLxLMwQ+Clt8Im7plaNZflAdeDE8FiLQa9u2yoqw2FXXAmAtttvks3heXmq92yJE
F1TlWifcHa7SHcIYdq88LId4ZjiPoDzRdcsYBQwGpTQnXcPXeeEHzb0C6bPsZrq88zQ7H0nCCGeD
NjGi3lAz5/q2CBRia8lcDQwAy4dDYGZDkmtJJvM4XZkVpmkMvoOq+PqqgMwFUTq8M4JkGsXpdnKL
KL440VN1P9RMkZ7fBNz9M+WiacRtyMiXXF0p39UwLyEUXbtBEN6pzb8YjEKOamT6j+MSe2yoyv5R
aPh0Ef+6qJ7WC9YQ1OkCSOmsiGrusZILyFBaiJ0iH0sTXmsvSiZ5Pc9V5+WaC+NY3ApZsditPssK
uofFHRgS4cQHukcHHGMOjLFLQ2H8i3Vpk8v8jwqMwoIsm7LCTdayh7yKFg7HUHUESVHjVdpYEKa3
5cJ3yeAhpNtyeirKxOU6hMZDTNb5c9tFd1O7Hhd/X9Gu+2f5mO7iHpYaRdaM65DEGWuZ+eOxXdoC
jqfZPkUP3aQDn9SKh0xUxv6iS1auvSTVfu5cOJEF++kucn6Z4xFZP74xCypCFzHHivmNzshm3XxH
xaWNYBnSuLfkoD+f/F58y44KWrQMKzIoYP4nQxiwTIXxBiYPhIyE3k9dkCuXMuy6vhVkemjuT5u5
SD6GOAtDBNvj43auHbKPchNtxyvKYVuOds37cqkDevQmoOTQb7WED2ygjcoOIDbzh0ymWrVJfg/k
E9MBCgCLEkL7uJYJ4ajyYt0fclsDqImRTA2NaoduAzthQlFnnNyss8tHrtptY0w2dSFImTHom7tF
x+na2TnIzWjeDTK5I26a+qcuf/OQi/8kp8O3KArSxNI46Wn8fzGCnR2x7m25x7YJ2JwonBYOqNio
HhCAwgeW3VJLth09UZB2ZXfg6ApZ+rXalLj9x5S+ErQDRU2ekvvTI3kkv/zCbiorVNEPJHGVMvix
4A13u5jYiFZibljgBxf/k3RRwzjZFc8X1hf7+lcakYdDi3Jv4O7MLl4Ru4nuV+BDVG82XWb6m2s5
ROOvEnKqmVFgWTkJ8M7A8ZHQHtIvd+4BnuG2Jo9IiQKJvqkaG6rcL/5sLpgRyiOHP9D98ZQ7U2uo
xBuyUcSq7yyAOY3C+/AdpKAUGYM/C4Av4SAXlJgWxv83rdLsKlVjaalxRVc2/sH6WYhpeAQY9fr8
dss/GTvK2VT++V8i/tJjUlLcrR7fzIVMY1oZsN9JaJre168WFpGlZxLit2jCvbcmE9fB3s2utvME
Ef11FzkolPPjxowMOLHdwETWT2hH+n8430sX12hkWwuRHpP/DuFGLeXHGU48ftkBD/k5hpv0O462
F7UTXBwllrBpjwYUf/CotEE2zWdUW1Dd//76hBRjtx1JS/WswXk/zYDMF/OlTO5ODkL6u84mZxbx
3h4HI5vBX1h05toyWdqct5K+F+rUfpICqvTbUzTFTkwi33qoERRj/5t0FL8UUCcJ905fMFHyECgZ
4sgcMHrl0bZEg0cLOHwrNG5UO5Ez9LraTTKHfGRPosuwGHNzVAUHKtmKaarw7WDr7zz1Km5TzIe9
kwyIqTB36qzFr6DzwEaOoBnQLtEtHqj1gpSs4eMpODw88mbBuPuYk9w5hIqSv6Cm6IiP7j36Mt/c
Buk6ky9glJ9aJQ+3U8b1XJnD20bFCRTZnQIJ6GDCia/EB0FTvgSKsmIyDCPHFT63Nw+dGW4dRq62
aoo5cFabc9mZRBMqmUS24FGDW8CurdmctQL2rydF5G7QlmJpzNFGItyI9EVdwHV/GvToKTyr4SkH
rhgyDt3/FG6H0vDaxq0o36KHSV/cBgizo89GpNnb3wi0gtIGEBIYLql0ojaZiDe0GC3R7O8bx3wI
4ojxegz4yjH65VwItvcNgZl5UZDrPJ3JGgKGrdk+cIHGYOpZavs1SAj6B/PT0H59pb2h2Sm1ZCCr
lhU+3lYUUAMTGgXtQe2IPj5Y1kzUzuNfTsl8xO1sc42FxHTyKQ84guWQzNkK7uzhj7JVQCvgnEV8
ZlYsnuSGOb+bXbWYphaBUXyks+wTxGGpl74yEcZpYlGFn5LqCrkSn3qjX3cdUFq8bHs7j6kRZ2aa
rwmOzq2u3U23DOE0tSVHaF0KURgFOR1exAWD5IBKFI+KgeAhbXdLq35hIWOLRTP1xp7kkve+QYN6
CmsoDb9SLAEfZydlOysXBGB8sWqqxMm+oRRUCgYrBBNGYOTZPlcfrcfHI2Ko7ggDHvUvtvw6du8M
Sx3ZAQd7eiE8blYX78KNPWVcFqrk5Fo8HHTQ0ycS4FmQhk5y1yIRBplZg7Z+/dw7ZYK0zoLt/x/K
VhpLte18tYmzmeRPjHqXAOKJ1oIfLeMBGRUMv98fdhj92hRuOsVhZ1cqdfMoq+6gon8zSva/1j33
aFCS7mKTM9Svp3OeHC92LxHm9WMT/P5NEOA/0lulO1xlHVVvYAuKxryIBRsWqm122EmLBP7Vcb1R
OYtB+svoAlIRWg7PsWiWMQFKgT1RQoAxdevg07mBW4LlPkUsXMsK/8FRlp9t7AbZpOqzGzs18WYJ
L11gikm8HkCxxXXhJKfYwvzFcGF+F2aOXdjpvBQK3/FS3ZtlP6pR0So4ejrX65NZDeQyOh+eaY/C
LrmE1mcHoaaQ64+fv2qile8hHUxnHUawNXbiZUfysZxD+r3KbApXuUkCD3ZK4T6Ca6+fOY3YnVYy
moAWgiMJXSpdOk0DP8uTsM92Igzz5yuJvV58eE9XIaPXyUG80GJGznWZJ45/9zGV0Gk3P1M1suy8
Sm7GrIdRciLp2a/hmo399PVIkfeTaQCbQMmkJUA1HWOf1N0pYfNhSAI3dUNI15TqOweN2IjRASlr
/0saGYqLQmww0Nl/0M6xJw1mPSZndF3sYz8FfimzqidQItIoglKyf1MErQFm0cVLA/7DWu9E42CO
eYlibfExWttO40qZiSVHbjeMJpP5PcrmmHoHV8JxDUG6xQIRIXqegawtKjtAkyo0KyNyHd0aDo3r
C+JurCiBU8twJlWimFN+8Q30YpqH3a6DhAXm5DiKkLJrwLKKOCd5hgGXYY8D2Qxh//i5X7P++iBG
ctsZOYERT+FMBXd0SCy3o8rjWKJ0DKgXtp76Y6utYqAuE4nhHu4n+vlOsYouSP1ekk5mm9gMlIjg
vsjaKyb9N0n4IGQy1He0tXa1GWzJJ92rilfqk6I1aoizu56mgJ6Fys4dDV39tGsQ0te+ib8UBulX
U58dF/nwk6YEyIBKNbSt3Ie47rn15dWy4lQM13l4cOO1Yaw/S+Icv7ZY5GTyijZcaS+VrjdpabbV
fR+LXXRFGvsvGLDpfJ2Pz/WnnBedVTb7R+D8pi3Eknz1cEcJkDjWsN4feJxTJh/l/1pTlXitdh1q
h84F1E3hFUMUoCnM/Z3O8/fMdtjLIHVt3Z1E2yZ2Z4RNYbwl4K49yvp7I5CZYjxFVJDvlwxH3J0o
BqRAOnml+273A9aW4sObzuiI09i8S4VQjCethPg049w8SfuXCEHMF3s5BB4BZe5pQCAVZbgfkt3j
2hX80YXC59rgRrqmAg4zn41p90aDGpYLaJwAa6vYfit5mcxZQDZG8Oeh7nX9of4EkDmWYtAXIsKF
hcJZ0GOI8iBdIe7K6t2sWDEV5jIP8A//Qo354Rgt3YsqQbPeXEEQc3gXqT550dapsifIn3VmtcvG
pNxy+YQYBgpte4m10PlXvPc3JzeM4rs6FACOeRe/tZvC+EjFAGcPqHFIzoKmmOFozV4JL6Q1iefI
w7h0ia0J7BcHddJLQY8p401Y+QtgzvacWHOvl+KYVGtrj0aS2jHGbAUPupU+YVbmNrMVtNbvG6PD
zOhEMdyA25jJZi9b6v1JAFPLj9lUZDGOdRY1Csb2WEkGIgWWXOfuu4UOzpNpw74Ji9hmhBs3zTTm
/82czTsBfTUrQuNzSUckGYNOrIgcAQmQO6WzfKIrA4lG7POZub7irFKgIsp9zPE2CwD+VTNyue5N
l1wguUasmZZBj8Aap63nGFTOJxe+OEJFVyjC6rrW1fRZtmdWb90XXj51BDv+Z20Hnu+0h1IS64I8
rCt8nHXXBiH+xLDGgvk1hPTJnpQF6p8Vyvon+Q3AIBX+g+ZwDJZLEdSJH94qdhlm6q+EPD558u/A
AuquH2hgJGGUgwhWhNmFjoIImX5Jj0F4WKA0wff/mdEpMBpLtclhaoQYHarJemD+Jr4CsYUsP7S+
x0gu0iwSlFNps3NTb7cD9/JJwEwjl/d3S9IsI7n2uoZmpfE8yJBQTMEk5eSL80FdFFiMw6bSNijH
wvw1AC4B0iC95FsmF6heem31tYeioXbej0TgL08/u5ff0Iu0fOaTkqsxHHECa6WLDNn7DcfvhRsP
aeSlMH55VL2n3whLuPrP9/HfkATzCTjAEC1W+mvidWGCmSxmDKvAWv4VOzHhC27KPx4LW80q0fgG
ulWWezvK+jp4qOrS3iTQo3E3bCmPxyc2rjpVMJX3AeQDONTd/hDMivi7hC2m3V68CD2I9v/VGnSq
Sl/4FDPI7ZlSGPLe+2vSBRdhg0sUPDLcbc+fKd9OJIr0qS0SzBdkd2zmOzvxgTm59YAKygplPatg
qmDSfp55rIsh2dbrdmifD6JebIBJKqAVMvAslIh1YSMzhTHYJD9raE5hp190TjdlEvRPqO7QqDzB
Hyug6yL/UTCjWaV1jXGqIwcvy5ItxgQZrpX/VAdo8nqTlgEZpyk9+pbK1Wy8+UU/0drSrRAUOVSK
AnmIg2/Ed30UWXAfEjGJWxBSSxZrS+GFELJuzi4J32i9xDcDH3ACYqxN+bXhIkU8NDtGrv19iQYl
cIaH13Vhi72rl0hQKNXneUV49HbKNMQfZ62s2P2/Y3L62j+f4wUgca93MbC+tqnVyiLVMXgUWwz1
HJTZ30PZRqrDogX/6rdVY1DoSQS5Pg5ALiInXJPF19zL82V/ZBt8177LpYYSC8g3kxdJvxhuVBU7
oBXWe4YClRK/sC6kFz9124rxEFba6eWkc3hlnkAh04wTtI4eBg8zFWXSob+9fFSGIg9Dhmo4CSoG
mSH4rB752fP3lH7+TWbXdnPqnjBrx3da3GgC8RDU79k1DgNlPwoaSdvPvNhiv7hHOjLoAUL7H/ZE
m6I4fKqtzXjdzjYJikV5flUA0YL9DFAy9gIthnqBqD+D1monhprmfmgKLW/4nSXsh9hQ4Kun2hkK
VC9ILLWI9mD8NVflWfC2kPPLGv7voVOgFbU1f+LqYAAWq8Kt9erQkM05pTo6aTOiXG6Q/0HM7T+2
sgfQIX+vymCHyISx2e5iM0EHtY1Bam4cniVJQkd213h0cZBssFaFAXZMYoEmT2mVHEoSg89dP5nE
TWAn1lvaavmu89F9dAlMlMOoWJz5X26l25sGGEq3SAIaBLRF2ov3A3zDou2OEfe9jVpcF78Vdv14
o90zb3TgDA71+rxg6emQ2SJdRnuv6I90y08WkMZcUVZ/U70PhAdzhIK6CyJEoJGGPAUxuHkAgSE3
eeA8vAV7Y0yv9npBzCReP0jRrRMT05+2LI7CdoXjC1K/0y8c2qaLY2dElvPy/k1wKtl5PNowc+Qf
RJtcrTck38r+CAWnANCh7fVdPA5inEMxMharjxdgZf7wOdsyPK0C7gITs6mcW/IdbD3pZzBykSS2
KkWBT7QHncrJH9ID45Uv+bZwE7I2k+aOmzk8Iy31zhCL8Cam+EE4A0WZLPlDHkILguJHK8Aiyf2d
4RllKXtSxXj/6DyTU29qXuNJmQvv6Jy7wWsP/XemvuxogCuKOUfp+C55igldTWzXp+BColi6wm9h
W58wDU+rGfWG5zT+orOODFuVQuhN/4h2kOtcK3U2SkU+XqoN/fiXqXnCNl4gDZHqT+7MzRiKbFzn
8o0I/MfNIkeRs/YPx1k0lbGoGX2EB3mpDStMZF3os4iHOZYNGl+WjKrh5HvNWS//Bp1QxNpJ3CfX
KmEQ03Ydd104aWHzjE+ImtB0tOiwki1IG6XNALuU5Y8524zHN/EEBqoRkZ1kpQ5/WNR4ZNXCGLg5
2QqLLSItI3Mwu2ewsIdpkKlG9YdJBWOWeeV5ccJ/7EVPZ6LN7sOvw9E57SfcMFVZSt0Rp0PkBQeW
1dpwC9HjIQMn6uH+GkuZnvNIV1it2grSbg+6DbnOwWAVlGAmswBPe7+/K6B62NVWVEDp6NRQsLNV
QdKn9NA06jOO9EToo2xt2lzm/Tucs2iXY+jwDgb47eMIkqRvbn5blUiwdR9cSS+LWRYbHT5nFpUK
uDywGAYUBB0RmCC4kCij1E5plHt/oeIYllgUeRRiOtCRue32Ndxl+0Ahr2lg4N8QV+tQkGi6rGZL
mKXUiA71JDBqasZpYG2CTYCoVurUlT6OZbv72rvkJ7pIDDN58XKz54wGKaTHpJT1Bc69QwBqp7MP
f+/yvx9GSyFEt2bCfsnXfD/yODwY6fHutVGPx/U/kkKJ2GYHq4Jw8T9uCDjK3NMibgb3V2JbcS+E
XWkF324eL7n07xBm/fMJdJ6sj2QZvbV+Qbgd8ShHe+37VNTyjOopgquaiVv2sC61Bhz4x/hKf2w5
IKnJpoXHzgAsn8E6PIHl1EJ7opt23k+uNOkVWlxMbBQM8HdiTKpfY3sDuep+OqFJ8pucfCuIoMkP
V0BtQq7T1W9Eq1/5w6TFTAlmk6PE8erTEmqK+n660O9vxpPbog+dQLIs7HpBk3n/UsIweNOTCxxk
Ue/IbUjdzTlYueJm/ANeDrYnZaKCSil26Ij6xQVjyLPYH0XLDF/zbpsygfWS7QcsA2YM7uDHtxsJ
ZD3hMnd2wbxH/59Z7JC0ATwVH9HhSc6QTsNsrhpSp+O89epKy8qQ2gHgZ6Zs4iGyfklseJC/QzT7
P/cPQoxy5D+Q6axcd4NK5hPurpIzlSFknp4z7SNmANpOenFIMI9XBJYugqSVhaqvsJ0DE4P8LlSP
qgBA9oqwwTsG5eS68FV8eeNhJu8OSlqq1GiB7z/Q59484ONjtmUGyUgsxXXQemN7PI/Bi9cPc0ue
wWbM+zPv96B9m50PtfS70Wo5BzH0iCPMamSxClXZEfCl+R4Mga7FKQgPRBFhrE/N9rEaJ9orHld7
Q8qGWEDhO90ysoVN64aKjE74Ov0xTu2MM2sXM2emLx1q6+F47iktsI5IU75Z6rSZjW8s4KM1hEIQ
IHQfR/T7jx6Uxy/5ZhxLmpkRDh/3nBe61C3z2QyrJk7Q7lC9qrs6Uu/xQ+pU3O73XF1KHzgT0Nlw
4jMPkeVHSN6oEzspOKrvtDmocUWw3k7vdL4YQcqzY5sgOluaJY4t85zIsroAGRWmKxnvRjcSiDtt
sTqmMKF/6pR/4ErBYoi12RV+KIcHmcIoT0pgLJ+4gk/SfBI/pZen1js0Kyqp7Gag3lnCF9Nt2KvK
hVVkkiml3s9IVz76OabRrHIKtAGaGPQh4KG8lxOH6A6rlnkYTLKLsiqUPVRRfbY9Ur7NitZIA9fY
cO8RjGxjMssWZTGQ0Ipyi6ARgLwnFx2fZN4360S2c+IMKOKV3Byn5vk+oyOZdNhQI3CbLyI9udUg
9TwQUgm1uMiqXgBLDxauoQHvBNRhLxpyJAXqmKut59s5CBXCulCPrLltE4Uk7iDFHnIJ0K4KJSBf
h4OiUuujVeawRb2Gm2ljWAZ8dWlHxPJM8bw86ENlJri0K/pRD8tZtP6NlS13144KoL2+agW5FnaM
RSIVB1ql3nWrYZnQvgrRY/in5xap9m3XYk8LY7r/mZmTtzH8PKedJbsC/gx1chZDSnMztuW2XY+3
2Wp0BtS+k0pEUPKlADM3tv3xk1qim7LR5NCHDQi3v1WpY6XAUCO+8iUggtKm25Zz1o7B+s04Og6A
BAPpt+5avTzgevOJvaHb5j1Wkd9fE5r++RJMZgRaRmKxgwjd8J6MZwprEKjl+q53DlDPDlytkv2Z
+KeB9GDKd7yA+/+1VnWTTyk6gRCDotfz30VUKLnIKZFliB22iYkgHmifJ3QhGtGcykgG+/vT9mgC
dQDg6djfIj4qi0RspDC+K7z0bpfBDEyCDE/Cl3hlVpykoRE10SeFTP8eC7bdBWR3Enqj3413vrfF
+CDpIGAhWdiU1TJoiJKN/twLbKPw9AqbE1uv76ZAa1HSf3Y6N62A4gjHeG0N7JZAMFf0AXHet4Q2
oYbCS3U1Im/+OOoIp7AN52NK50Gs96LXgtzxeLjl+HqcEe4JRnZoIu+mnXgp/GMMSgEm/PI89Zfd
oN+YM4uRFYDMzuOJn6aTGHjACZ/CuNhwCsc/rg+uSy7wjCVhN9bDL+cuuYR/E2nguCSUNN4yKqp8
wEg4fjjwMoIXwE4YffjSX7SdiIxbOTkKLdQV6m2MjQfJIkb+LLnAdJ2DiwtiQR3IKZAz0RoA+CNg
zv9kB04LX6OzejiOkza6pWL42IKyZjgvyBcn7T2i8LUJ/EeYi9T0p3KGbwUjE5inZcq/JhdoO9ro
vsUy19Qfr7BgG5rLJ/p6CozPtMOTXj0vlI+G/VpPZL84S/OhNWo/wtKO5EG3+XQ+3pLDaxsG3vxF
FQOVolpd4BNLb1vTqJbGv5CBxZS0AcMjGqUIRY1rVhEqqIPYJfLP3kFmJzqLCtq9/MT3HbxIai2I
zBJb2qln6t+/bZNVHJ7/iJe9tj3btm3Lk9KBkbGsnx9dTQLnBenQNyHvvDSaF2+KMWJrRHoZkP3E
LHroGCfZpGQ5pD2F8jP3lCvuADV3ZydbSoWrW8EdR+k7ygLKAEdraYS7Zied0jyf4MdEJ7wMARuK
uYbKOazvM52Icclq/v/Ce1yp2J5QotF0huwd7JqOuuDySIISQ5+hjCX4x6rkMtvVTyRwTtn5Yv1Y
MH0yBlNJirDfYojHxs+fWM4b3leZARtwBvRbzHuGQ2waQgEICIkb7PEURSn3wTqhjBnosLOugiKi
Jq8eQgYAWVszouMv638aDkYuZdOSEZ2Q6SnGK1jFnSHwZnBdgonFNWHR9uZ9I9SeZ9sjawW5q7PX
Lb3ajiQsVaPafxP9J/ud3Ad/zxOeA6sQkFg4ARBgmXcnSwEitan3ccJUkPImMI2KdX8PiSSPU2bw
NgAUpZGtMCpT9hk8jl1CEk2Ob7YlJ7FDjn9z1wj4BsQ0a8cuitUE7mkcaMlsQtFdNYNUXG+2eSpU
T+9ezgyBqijw70DKdd9+NtN1Eqpf+ahVDIl+84KHIVXRdJUPQsACKmi0TrGHFDHy/50RrY0QtclH
sjoiu2KdNXtu8narw+wKaofy0F/NV36wkZQsmyac5B3wNbUWfM2F6FpU+xbrwHGkK00tjMKgjnZX
eaexenFLY9Y0RkbxJA3wBiYx9ZbPg3UCvac7xzHtKYUzkEGZVd+0k6SEZjk+RD+Jeu3/JRfhosQ4
p4BsiAnnr7OgMNXawn1c8P1Y6Wj0UaWjJ4a5yIclMD03JVOht6g2mWBKKg9GNfSTHbw9ysXtUt6k
aNHL2bZr8/AaRPd5S495ji3cysh2/JDKd+nrzpFD7qKErHU2gs+nFx91SDI+/YdLOJ7/rT4mLIoZ
Xphddmeqb8gyO8qRYyOx0kaZD85nZdq5WPClVeY4gHhyF4JZ25LWj2xZXkRuy8GaGCp7rgnxLJ0o
blokkn4ijuMjOYlizEX+tuHsB5VmITKcNw+2ucfD+5/cW1Epzk0p/dQDvtbiHpmAtMadTQ5AU0Xc
xZTbMdMGjpNwBW+UJHam8mzyeBuqKpSxOpeAWAR3ldUQc+hw2juCvZKCyO9DadqyofXgXrYGY5p5
rLe2vlSPsDl82Y35zY87BrbK32GQTS4kIf5u6lF/6kpPLKfXtWuTskTkl7ffx39Lg3rBHx0BHcBy
jOvEDrPP5JGKc0TGLy5vk8GRK7FoGpbyKkxqXOAI0qTErFUV+j41EynMSI5UV9pX4pJb5ZGbgCu0
+N1yTQJRURs1W3cNkE9XBc1bkC2SLBAFCWm4FX9ZaRPMwJ4ZQjXseV9eqSdlL0Poe7chcEEXq2Bh
mqscxvK4W2ZKZFHP04LRxtlwYcfEARoHoJjMceKsZyUAaQ7caNIV2utLxg58ou6BtYtO5PCnM/uk
xozRMf1CL3HEnXhKaaOvMdhLVXu6WMj2CuHzmhJoWB+/1ijxTngTAaFB7NY9VtDQpGAM3X4FHuHv
pvLjCjStCZvYuiGYlOdYTzDaGWNNI0rTY9JgRg0BkpRkDMHHJWQVnIXlMv1abrH518Pt/eOCowG2
k9Wp+m7gohP/JTMy5idn5vwGdWZsSqyV6s7PHTCIAeIKNpfpxG6fcV0P4OSyBJG4vXci+Z2gAqkA
kh3DO6HGWemUQ2XGybKeveZ1IpRupAzoD9XkOgKvoZvnzylRQE/x1hG4foTmKyzIEFWgcdmaq7zM
X79YOHZ+B7y3H/rs0D4OxpKBdHUodoVDlnrgLSX+TQ/9kgnbjRfmtbIt4p6WU4aeSSzTXvmKNWZM
924gMOxBEz80I8Bh0Fr4HAccPkn0fGXqC/oVNHC2HwqKkWrIGu5muaJIhwrjVoJG4u7qAqJepFBf
Y+movfWfwZk3lfCKUU7tqzuqu+x+eB3lvqlE/piHkyspWPxdZ1qIKKKOKltWCtRbKOPuX9PO6nFK
k5GdW8ODJ1QLDsrZbSMeTVrn/IHaB/S+jz3opy3iTEmbxKCUWOiRdKQ3zao2yKIJs7Xw7gIjoCCz
IxaEbjkeswpxQ4G346ZuAjQPuFquF4wiqJNbG58p4tGA3GeF5/B3RsssiiGDE6eKi87vtKR2x8Nw
iRrn9o6ypWlY8smKjjI6oZ0l4Xt2U6+/SMgiM2jboHB75DjsA+R03BkdqmcJA1bCoY9ENzPcG5+/
W9+7P2O6eESnvSCh6owDXxFPBDPpNEcun19jqfyTo2TTpCOGloU+B39/tC7Ob+w+zPMg6Cqg03nl
tgvhk86f1ehjV3pQIOfr2QbXoS4NmfUF+zxVFtYuOSo/UqE6b7q84XlY0XHgSaICYP+cM0XAiAl3
L5HxwWF8Lfc5sYXnmOChCRMZ/dtnPiubOCk9fr7QsQnBB8n2hGw0031Xpjc4nc/HUdJK1u9n7s5b
FOvu8FIeQRLMdtGcc846AJ2OqRcB242HbGIi7an1YR6wxZp6AU+ZGUMLvyqLmWbsyJQitoOTnLAb
1oD45yCgkD+rL2CkkW64wdyMBwNNAQVP6LFohD27RZr+RV0o4aFUKENovGb1CVyRK52oWtE6HNb5
xF/Ho/31Waz0MkKTSiTJo/Ie0vdUipg9DcuLpYGWOXytApA9s/aojp0VourTygt6p/DYUDfoEb5z
j75bPalFEHyD2VbcB4r7PPtxk57pOsfMKiZp8ksYBw0q9zzW9b9GbS0RUUrIHsui1U6HimaJoxj3
7BVwDovYzYPsXch2nXWacfaIj37ET6sVD7pQF4dUttwT+JIGC6pG+3Np2BRpBfstPlqnx/s8gVFv
C3tcwHTFz6MWps8AgABMO6sSI3c7NjRawq8F7WTwoxQ4ym5XJ88+vjq3TRd52Gi5IyiGPgSisTxW
LG0ttf6/iw1vAPn4jOiD+dHCfVk62L3uWYSXcbeGs0mdiAaZI5MChZ+HMpR1ya2TeJTKakw0OUcx
twcyk4jS60vYX5rdfcu/uU7Qxh6WZCT0H38L8ZYS4C9AFL3/yZsMGrJxz0OB+keg59LZg5lnECXY
XC1M5DkGrwa0sDZKUjPVD4eLNZjtSrrPdVRWiPz5me/2fvGa3bTdP/gsMI+SPYX9iWtM+pLyHgus
8p14ZDAAKLFyoCKCLssmbHtPOshtoZvGK/YN9XW4Hh9y9+IByNjlTuw+b1fjnolr15iU7u0B7L6z
/mYQmG+oxztfvh8A/W9gSP1UZywfFB9IdUQQMyvCJBQLeBGdhONq4HEOzIfYZ/2Ms8RpRBJ8qROd
N+Hr35IEMBPTwultvWRcRRFa59Yc5YEcFOIXNesbuYP8FqAF1Jhb3KJm8+0jO5bNQJgv0zjPE4EE
6bLtoUWympKiqP/Nc/0L9aDIqELDBIUfhHi/spdvT1GaHY5qA5Gtcc5YSkce/dia9G9o7xDq17TU
1uXQtWdQc0EsoSE6aTcwLHNES1Unpoc4lVDQ4qkkMXh36ltZ2vPdedlE+a1Bo72PEoTXLAiuunRc
bne59X/K83QuFLk0Q5GjFruzUqADkQjFArDki2icseB5YMhMV+CKLKEK+VbLy/m5biEgHbuDMTIB
EC5gdfLtO3+QgokJRPgN3657Yi0sSTcqCDAdbM4gNm0CwNXxnM8ycSUzasDMW2IAW7umaWNdhbpo
YvKGJYkZptUVdf8zo/uUTv66mxggI/xjQMu4sAtveWbooEYS06e7yTrk+E/IIBhktKw02mWjFWSE
EZ9adkb8kcBOBix7mdMjTqf1a2uDScZKTMvhDyzYEjD+OjUPP9URL/7jU5CdbBxYTf7S9Fck7Eli
4YxzxBoupVIfKRXfd4n8jQ0U99CqW6sN21dOE7D9O1PeuPALxMEVayGZ+aQRDEwdQr8lRQZNycAD
oayxDyIL14p1XLU66ROkMoor/qxV7bqWandkGYx2DD1j5ZTYs89GJWbVFZjAGYA1V+/28kZ+XE3I
dCTb19sfqSAZO99AEKD6/lsXh0BXb4NZP2WFuSnPCIX3p1jJxwP0RXT8+AD+lddohiI9KIul5ZUj
iOhFPYfMV/1xE4ryPFxmRDgEs/bkCSZaRAXuAbpwhNI4mCilMImFg0on+nV1GXXVGroGLALkzTlm
Uwk9NCQZcJhwXThU0YW3glKw5vbrpnVlJ0b1WsvwMSxzcAhIkbpjckEP6PNRLjSBprXqSgrRKBOo
3XPPU9uGrL6bPE+2i5LE5RxdLUUJjztMq1BC8K+Zo/Vqi6yJysw66dGPivWGZPMCWzNPtOhcJKaR
qX7GK80m128ODk/xRBjcph1bnVgSIDzuWZwcZmykxg+VewIVHer9dIej9ih8sQ1EXRlaUIwfjP+o
0xxsFBJzMICHWBvS6VE45XF5NV8AwORwK5mQbOoIHzpFlfQBVivFbP3U7ESzUs4YKPPyXksBnPPL
Xx+eNu6kxkOYt+QMMC9qKQLFWWWJT85269bRWBmL8aVGXbeeTXzKsW4z7ZKP8vJ23fJltWFfR26S
KAZNQxRODbZql+UDAaHyhPUP0MW8aIQ4Zxq0GfYqbAGVTc6E/pJojwvM0lwfxl8HXmMUIW+nfGNi
ZxQuVQI9D/qER82oera5KQ8FQ5zU3MEnwGsPmqGkg3ZufH+K2vpb+oXTiK9GNZ6GgTtBFGW78nqe
4HRP3BkqOHVbyVwDOcyBze3sB6zBdhtqb8+4y4DeI2rouJ+OPq4ABG0305x9VG1KM6QJaB3VBGyQ
5nuXat5GZ+dHWzwjdYtOl4dVFGESmuPoYSqvxwI4b5TM/TIPO3tSyWFAKYQK4rZXo7wvGO5lBqad
/YDlaUPuYzTDOld24T7IAJdgIxJCQXopDP6gcnVjE3x+G0f/b1gznmatavSNzu2vvGL2tLeh+WCc
HzvpZ5LGTHSA823UcFtaZXMKH+NYoB6ppyqaa19IfROc+zHovKQvrPCk7enxldR1Rln74f/eBD5F
VvU2DgX8HDhSDVZXTu5KcBTdZwArNZLk0yUgaZRUyD9yf8kNn1Uoyb1WDe40zw7ewdUkIrYbteQI
xoNb785mJsnlDbDd+Gi+IonmrLP25B5EkAbD5nLUs8hTQEPHDqZU316yMbld81Jij8OfeqjV1t1Q
cn2H2j8BRJZVFRjXSN0Jb8P4zZyCxh2i3juSSlY9kPM6wPryGLi3SyaLkWy89rzdmrHOzr1oO+u3
TXjFQoJa4LVye0pr+9PGvCQD1PbnEsrUy2mlwHpUktCqMUpo07kdV13iABzZZ6ybUbSs8waj+Hjk
UFdJhKdcaox+5/bak8naHgvYAckcvLzLnVZKi0ULHJgPQ4IqHAY36GWkElTiYkW37AMtVVkL2aoF
cRSfeD8HRpE0jaDpMrd/lkId/znuFrcmgz3dNLWweCRJ7JkNiLfsFMX2ljuhAiIms9Lbwa0qPC1I
rpIcRaiE9vGvz4sWpIPpFg1Wf0h2ekufNCOgWpRYj4VoER8kl+rJQh/cz9pF+n8ue5A29EPVjLiC
N9EvnJKfggDZGXWCm/kqSZbGv8GS+/v5LvnCIIJ9TZu1SIMinpBCzlDZHyGf3cRy1MlBWfXuv4sx
+IgJoferLP72cPLGySBxgyBwaFCbIR0PxNZlzM0KZ7NCCrSWCiVExUbYcQXvQmjxkamumNOkYJ37
TneTs+JR5910BJTrob3kxs/S4nof51GwPGtI04Q7fLBKuZpq3eBFKK/GokdyrrWg5BiAPBecx3h7
og4fZ1HZRJKq0ImaLLLRc7u8IuES8rPGuPOLHCXpdXJoneHHxyXEmZNti2JmrhCjNWYVyV+9BEE+
nZu+MAQ7o33JT5Gn2xgRboMfWaDyl/1TFwXFs/1QgCLswGNL5n8lJrGL3DHqqBEujyuuHFasPkWq
45it9WsgaWvfG+n5Wlc9v8O+5nKFEU9u7oAchhUNBDPvOmHi3EqOXjgwbs1dVRGLqzONFLJjqQ+r
L79iipO0j3NDDQeUXPiZNV3Cd85Iilwfn47378Y5a8++FYwSoivcroq9o8fLzhx5yCzaW5wOzeDp
L4R/WdOgvETkWlDu60gMd5BcxOccxIRKGiAekTxwB4RMcCVEpVt63EkoN0GdOBhRf0R+zCvjnxRV
haecxeyRABdAVrlgqj/qKdTSXP3rk40PsftAEXTHf2n/Ir9VmbDJY0JfIy+k1sc1tnxEQb1ujExe
wXV2rqp9N4I2q3dMaHzxbW2DulrSNdnXjdZwEPDD3ZRS49dy5wq+USIW3BAA7xmiF4VE5mkJddO2
6fGygSFVZk2KOeBV2jQJvQjidmzp641qC7QUq5rzimVhjajgDRH63qza6JjB1cZlODlHPw//84qM
qJYjrk3+rPf1EqS7espcpXDHEvgX7hJ2Kfu49F8SqRSx26FHgUCYDBadK+p6lakVxq4ZddsySb6J
59ug3/mZuH0pQSp76eMFmsNj8HgL6CouRsHmViQwSp6g05pdaVe4EfqibSiuuCbPG5rMlrmmfldF
uRSiE/dfR9iSkJsKz9eEe6QBAQxnf/78Vgh8GciJwCEbdtYVvU6ISuBnm3ZQWbkAs4jdU4FRfBXl
sUURpSHYG+VRvWqae1nh4u32AstDTfVd/fYu+OeVcbaiZGqlzek+IyUq0lGrqZaKhfP9672BqRYS
tw6PZuonWj1nxgGYorsGgPcYC3TN1/IzcKgx06sjkDzv5yUBgVxRCYY3W32ZFddvI/BdIR28JaMa
9w509bTtTRftp0uD1fYuBq5IyKzf4PntimAvkZaSptlO6BKjRXHVZQyUeaYsJse9wYJO9+fz+rF9
Y4An38Kmf7SnkV4wTujwO86M0gz+bpmSRfPa5wKIQDfaXDt5mrGn8bAGbGOix7lp1VkX94C9Vool
FZlR24/Gj3R74rfPvSu04F1w6DjMA8s59wG7nNLfJnaWIHFAc1Q+R0YHx0WxGMVd+LwmNy9ytkaG
9EPPvKcuFVix9aKh3aojRErcZHTjdmFa8Jn5pahz1/JR33BGN5Vo1Sm6RLMVsMddi08RclZA1tz7
UTFitgsoPctetiLAieevfeBnCkiKE3fStyuWVWNfBEb0yU5llxDvf1NkvT0knHgEq15uH9luzgVi
H/AgdunGpxxnlTck/RkQtki/XUodYTF4klV65aeecOKNU+PHa9/j4bfTJfC2aAtiMJP0BciISbpD
FmM3FJgc08ngABlB8Y1IB5GulI6ylEYzsOyXX4qlnt/nrLntbfdUb/JQ62JWGBlLaJZ785KdtenN
I/N8CVu+WCJAoeHPEogqIQnK0QDOYs6o6sVy4YFnNUkB2nbR5aoeKPcV0BLLHo9hytqg3pJoosY9
ksOeI7mBcJKZSNAiWf9bJl5tTL9q5hiyYaNopPC8fp6nxy9kWQV4LAqzXW3FO9Vp4Wh6fJUSE3Pv
mV0to7O9NLtiVMaDcBd9sCgKikxEoyAoJMc/3y5cYEO9TKOhv0tCuV4GGzdQPSSe4wHSdmxDZGm1
itdzssun7CEUBnCj+B3oPZ7aBOYeD3M+bG5Q2KmUNEPRyGOwKuMi0bi8hHBQ2BsBAEZW7BJlunRA
5aH5sEtiSBMYndq3mvh1FgQnqKi/Ua7F2Q0OmS2TxUNRUpF3mR+ZUUqnvpYjNBM1mbZqCGRT9hdB
micRw6IiL5AhnxuBUF5eMtgvwQaAmFuaP4aml8wW0TxfimNuqAFGtL1wyxvu0656o4swGMb8pomE
sPF2H+daMQYqTiNnq/kAzPrlD2G52qj9pEazAANuP2GOMfzcQPKsirxrZz992P7sNIb6ScykJmPA
YTab14jFDEn1TeCPLWtH+ZuBQEMjILgLundH4wffhkBGW/69b8+WK+9+gQWihnwSVvSQeiXVx9AZ
0lpEjCii6ZEI20bamEY+mEDc5Zo8frcP9P8DeWYazGSw+kockBS6uFUjru2Nior7rOULyOSBxVTX
chaSbb7y7b8+O5CUheRIYShpC9lH62OZtZuZIRYq5XvmVOlFmMlqgofyBqfMRMQVsHagb3EiBgOH
mQPYLHN0gCQcXKEoqMAHGLrDqa2Q8G+g0SyksM+IcZ6DX5bgwPvihuoJ7INQMvrqrJLflF7BsGuP
HtBRbUTSWYusaICZ6V/UWSvdbRjnc1lQrN7b8OQi1/D4IcZUkIbZjEPftMsQNCetORJRkMjEJTCo
mpZrCb3s4oOVnB8X0kk6UnP5U0s+qZNOTyqySMZmSdfyPRPaCMOAME1EfHLbCHyur5aWt7nWc7sH
x/qhvBvohhM07RVwf4m9GdWH6VwIzsUGBhh49BbDYCXvkDzG86ntEtBLjaSGyfF7xMLyNU7kVXPO
+D7FoJfwr0WHnN3YgkKEZRsGuGwOn9ei8GqiM68bv9neohzMhc50REWEmXqB9YJI80ig4ytm1B/L
13uDdxHDbARXo/6E2/vd4z1fNJsLkkneUmOv6ujpHhSCXEOBWQK5n8/JGocTjKZKozjMP0tCV0E+
stBWL0twiWKp7ZZ+njFk6XwC0UCxBq65+O9PggbgDOMltOwML+yw6mWsPfPAnRxrZY5G4t3mYq5p
jfs53OpCYky1giZgL8mBecr9Jdp3MVZz08VM6w0zir0LEbl7Wh3nEg84YN2nLaiYvL+fn7qS8zP1
3v+LWPkCAZFqKnWot6bQfwZwiVuqW6ej9TxQ/9JbpiTedUpVsAE1P3oJiPbh/udDRr71jgZLCXvq
QPSJ9Met/AisFbY9VMAo2zBFq6iinVZ+cu5eQkuzKW4GXh+sl5XezdyEzktELJZd8ODtUmKvWUST
WDyfE6rTEr2hkzobT248/BtVjwRp1Qy+IJ+/VslFefUextdextbuctY+ZnHLZjGGMnuHa8udQhjB
r8oJQtC90cFSb0w6jzuScJ7LXZOXk5nC0L8U8CS4rlJGWaTmKda28iPKhV0dZaNdKqNXlr2JFkAZ
gT9TT+Imt4jK4ad+OVGdagQpLGpvtSha4JbMQBmdv9VOPksa4s2HIdb5d1LZX1XsXw8xbHb/3uk5
hfwpIRkbveXNU98j/S2bFxcs3R53xqguc1YU1Cg9eI+VktOt4TG2E6EqGEUa1jsqHxeGULhqFoJV
+O9gu34VD4sUe6/fDZkwYcliwnttUE6nPZIobBemiMlCiMltZua3ecfw04tlEsMguJnQzLnZKPUz
JaIRfPlFJ/nKxjwogdsTK00EEPVJvHEV014hU2Hxvn4hOeJyWhpIurxxkEJqdVCNDiLCPDzTqKG0
JbqBeVG2/qFIYXQWLdrXJvU+TjHwx5FNECfapbqxC9lz2GILtrQA4iNYynjpjQmDWZJKSmssB9ZK
UxiVwn9uYqIEhdpsPTuejUrV0pS4uLAZkYB2pufuVJSmOJ+Yqf8GEcuSCaOKY8tl+zgdmJanaTo6
Si8vS0AR81eSq61XL2sThdVnLAWcqEr4Z+nJhagH/uzEAMHQMYgVTIGpqJZiWXHEtzue4yFDlhlv
NKQmMde/x4PhMwdy6OGVzjOo35uFOBxklx7TA1qpcOXU/BcSW1sudgWPjLIGE57ifTaYHajwVtBe
3zHbnL3rgYAuNs2TUTRinuARVJldH1Nu5Zi6TXdWS2fHfwGNae9UHET21vjZgQ5AnurXYhqmPT9A
CQBFuWc+iW3QIN3dtwxBHFZVpx22JxqsS494YfVFEJwnc8xC/T0vraFh0I6C46bFWm47R7sDG1KX
8MgY4g7oqW7rsSbOchOrprneMI4BpiqBQONgJkMGHdeBWDNmIvZYmM+A5nDHb+oZ97JLTgIRiA0Z
ZrJVQ2MtHnfEYxCidxY3LLL0u2MUDSTdAoDiAkIF+4/1VTOvxz94n0M4m1Nw6j83wzb3Zd1R1E3D
7wLiSu95KWwQ64HYujq2ndDDy2LL5IkHz5//+X1fYL3Bnm8Tq02MGCNOfLQ2TaBsihuH9eVJ6mar
pyG3H5D6xyTFItEhFsUUngvFwRKcBON3wGO+g6X0cAt+Jl0KdHc9QqrCr5fErtCYAHuY8Og5oGQv
ohT6UwLyMkeLyo4dwg+WB1T6vf7B8LIrwWLBfBNIA2dsdd9ro3GT/uDX9n6jP+yjTE3mUQIqecQp
wl80BFRUnuIPhJrB6k+3rp46jCAWh9V680PtORJgvMd8WchRoDHnESq+G5u86ggwYSnlGI2Nh3wQ
VsXMQzjgpeedYDrHhlTSd+VQFCyqyQcJL6bSTDNC6TkD14KUcJkpVpseN10sr/ovYaqMGyyXAteJ
rU12uc7wC7DlJxLcIuOTPSAQRYF87+AgLbr0K1RPO1/6m0UNZLKNoOaooclb0rdNcSCf6fqxVYxX
T1VjTAY7BN2d+qwKEOCbrvGI/fmW4WEUR/GzKCuplD+r/HXkxKac6B/J3OpV5fhCnPI5pd4kcLRP
IeB7IjQDkuwVjDw0v/wWeokwuOOwEJux/8zo/C+SflqbYXq+Q/m8Fp68/vm/AoAi6dgNT5sIdPMt
lihW0O5qNbqkdT1d1d7GZLi50w9Y8a2IdfAQHEWHx0gLKIS2dLtIfu24EFZbjBoHeKOpG0m0qKDH
8GP2Uc4qTpfdFw1j/MXIgWTc/bfIiO3Ap+76w6oJMwpL9BW7RDGDuAsKARAEzPtMVEBYVpIuvuHU
2uLza4oEBOs3O2ZPQVyERdR+dI8qxMUhy8NPJ6v5Gen5znh9QVxsM3/HSmgBW+Z5u2P0DRi4JgbE
y6KiQUQQkX+fTEbcxupkVzQWSN474djd4Fss1hFN9a8t7cfH/08/MSvw7AZvnFxqVqK2lZYAZSku
XY2AHeF7kGk5ixCyssyAXS+rdnXY4HiMNFMCJyEElYSZESfWu+EHdBwvd7MlYZeHBmqmHXJFWfo5
fsX3zQH1CEEZ5t00vHE+zIg2/JNP05aZ9AzbSvvlu6ja33l52gTdtc9vGLs+HrVubkitL/GbIg+8
Uwgl0RIwSB2WdTupRcy8wulPg+wo0lDQe1WLSNQTnHsfUxv/kxh4+GyOokUqVKk7BwQ9bKXi8HM5
xhSsp+i1nv9qecJiptkttkT0H8tCPy+scmE8Ly3NsQKnLbBTOKLuG1LjiZmz9kExS70m6hYHnyfL
l3IDK2KqPpMgClDozBIkGyLF3juFZftsxBQMYF+41bDZ4Ad4ATx/9v6WQ/t83kwXNlKATjweyKdB
GI1PHwiuid6nFwK8zMAYx5PmWQODD0CN9ZmWNX5jxu64DENdnR+mlM0f8MOeHIJTLaI4kz2jjiET
1/u754VYmY4XQ1NHtKL8FC8pTvHsVM5/VuTOaukXK32jf0+7MCJpSfPWgDu7rZ6QsG2grof6XIin
ttraD/hPnefgpy1IgYKCgUGd4+m6s8gk6QFSrV66CfbvWLV97HQbQ78Fzsy/a1kmlW9W0m30Aqmm
7+dzxZ6Pgrzr4adDOny5dQycztPPsswRTMQCf92AZMls5f1abc3j0gGzHdFICk+RjENOQWW0UzHE
XhecMb2Ubo36v6rT/qg5ZaeCZM8YfVg0WA/f1UeqF3kFgcOUix+k8Qu04uKiJphsK70fbWUNXLtH
Wjgk1lSnwslxlNp9cx1Mb9bapBlJoBHVH/QA9rUooRc0Vx4gc31tz1KMdSRSVu2dG5nLNA0vP4mK
nfzO8Sq1azeBCmulFtminDj6zCYBM1Doapzx8cUifMaLgppsxGr1B/kc7jO+n7qv4ee2CTKSB6TD
bTX5t+tgR2Cpywg8sTOK8Be15prdUCilfOgt94UU1/fUZKCfs2sI86rTkBUsD0NmlS+8mhiW5voG
PzvV2Q3aWJS/cQxicUX/zkhjQzWN1XxWAwsUI04oSidZnaZAL5KpPcex2NxfV6CgmvSaT3rhf2ea
arO9P4UQlrm0DSR0i3rBQ/rF0QUirvJhDW8J/cRvlhWIrDO5LlcEqttJbDUGXe5pttn+rCG+hIal
36WIPinsgDgw1Y9xWTrn8hx86cEAuTfE3o9s+c3J2QlHQ8s9LLxveLyXW82pGNrPGhaq1Lb6ySkG
0Bx9fRnmhyAZ39S1ykUNY2NuZK1NEH98utY4lKnqKyCdoSKvvV38UhaysINSfSIIY79T+vBzl5PW
gGVytjAm43z+p8Wq4hFwU9+0YbaBDiAlb0JajWiuyAlvU92WnbWy7d3SY2JH6outTYv6GJgKTdFm
9qO4TVxvfEm10TM2mf+j0bZXk1CmSGrYzN2Ud+//h464+hjehNwQxQTsvg3cNlobYoCITiEbtFVV
RJZPjb6vbTKM1IJWWgCi3MM4ALc+7VQzJPvrq9PCELfR6A6pvcX65oyq1Ms/TSLmj2kNnGwMllIx
MGrCFmBwmmTQ9i0qGA2JqdU8+A7625MKdRkcXhHmttCoaeaJuO7Jry6n+NjY7g1WPteu0C/X1Dcc
Uxr321ktOti4focXOnm8mVQjsGbnhvtcdkvAI/RLZOZehvPAWNw/mc3MvamaxjkT0NyDaBIFzLL/
ciaBc6vUKvr6WkYWrA99qoQ5hAPTeN3aqbGMJ6xBdN+xEkL3gxur9sgOTO2XA3uxwJkw/ino36vE
uUlgmPACVZD63mw4UG/mSTe6dTu2aBI4urQR17sgyDB7+euRF4xsE3hyGNK84jSKr+dNGRP1tAex
NdeMmfaUeb0mWNeGwdXZCGrnd/Kghz7DAFmtjN2PNgJzsXGzJZxUegh/Uh3GT2UA8KSjXoOH49VG
dL54ysHz0szAinO9+xLUuk9IC0niwzZojsj7qAK2L5LEuVV2/mqUYpqCpnCTzQ8PU9cOthG8bXYt
/OqPsj3NsAa4dGkkd/6Wgk2dM6aItyHd3vPBsqM/KBEh8euBvwg8JaBEFEpp5n2Jb6nY0tFzj4gV
WK7Vj8CdZPiKcCb0eLTHd9eZszEoiz/4g8NvnJoqqbggHg7HJPthsuAVJwCVQJG9vG8EAXABfdfp
4gQUMjhDLCAJ20hWbzEyfZlFbSGGXi8OzUofEgdjdruuYeN0uXi5VgHgbRfz1EYNfQUsS/3DtTz4
tlITnFZBl51r01AHLQM+KX1oQF1GeAGPxejnKiEUMn13Wqsnt41FqPTqCaH3FTZnRv2hTAhft47h
OKs+gIo1LsA4iv1lodSuHumG0Elw2Ru8xCgoSa/H/TgzAt63PI2vVkxlSxzl+1t7M43pVlzczQv1
XUMY6xe+SXSFvS9aKs516+CSotSndQA8zBh+YDyWdysFTZD8RFx6cxV9mnEU77jKcnkTMVmxK6h5
xIhVjrqZ2x+zXnEDlLrhnEztkfshmEQs+Z4fwn4uKzPBhF9ke6QSoW5Fu7PrlGbSAvCx4wyZGyQD
X7iR4Xo2+5R6JDHTnKq6aIrO1sGJrcpp19Rr8z3+qZiMhUHYJuGyzqdEwwvz4ISu4UeWDdmMtwsE
1+w/IyFL+hbIGEBf7G8wPhOn6e/Tq8zLU32rfbiqirfB2G+X/PY2GJvz14XW8tXOUofEi8IbMvJF
+FxoXPsjm+u9S4yyRjfpnxfq9nmeHS/Ck3MGPPqZnM5pUZUa6407ed+F/WMP5jBTOkYY9AZo/mnc
MHONcxRumpin4nrLccb5LgHS3BDHQZ7tP2AuNuTpOUCcaAqeN6m9iPbmddd1THirDiXp/7wKdk4x
HEBDoJKsleZc0o4EqwsPg/TZoEnXN3NOZnJmtC/5XNqzdQbkxExkmjWhxCypu/KGZy0/Gt8+3oiN
WEylK0izHArvMMgRDny4aLbnIdn2JXopDjyeW1wqWIW5qlOaX8pn08STmxNNPF6DByg/moRGFJJp
58Vss1Jyp1SBTqwqJA/E7lsF1qjVHPq2HYjCCPcThTh5RT4mq2wRkaWet8A4IfXPcAGew/mAQVEf
0XMjZ0DPI8HjuzPGlxuqTj/Z+Qzc91mzcEzJyGwzVYr11/a3y73NOisC+ZTMX9iQqvukG3Ivab+f
IKrPVQlECb6KiCjKHMKRz6laDfV6Tz9wrxaD/BHYhQF9wFmL1iPDFRPr3q0qbmvWcfLX3C4+leeN
BZWfbRq5N2IzhSR0lMKZ0MhDgxN9n1kkx6Ssp31kmm5FowxH/J8+EHvA22pUlL7ZYSPjjHaVYH8W
pKaKa5grV5QLx7uQ7n3fY0P9Nk6WuWw4/3UHC6BcRR2oiARaL3gWc0QQsgTaiLUmEr1hR0j2Cbuc
AXn4OsNkfdjhCFr33n+TzTcCIOYLCD4D6XBHvws9liVdU0zBOKWyupK1Whu9JBul7pzapC0iE45C
qJqVCiIM5/l5toqB34NMMHjDSWKpcfCo59JEPJBI65PWhk47AKhxm+s21aEYnOmpLFHGCrRR5HWa
DLuxEE18qH/0e2Nikc2I7i5wDfnT5bgw6WrvxlB5C10QJVkS6FF1KHoGzI5DAwwY5drF4+Zlw63U
fcPTZoffUsFeCGvjZZd06TcvxZf3bscsuKA2LWih2XbcOWrLCV2PDiRL6Zk59jB/mb9xRVggeGE0
RYdqa+bxj81EQZn/4R8qCooUe4a6Z+8y20vtQ2VLf7kQQ+l7uhz7LjkLOc0O9MKGrZ77qivNWayy
Vx9+vcEBne4iy07WDZEba8qBYaCxMlYgAH9X4MI2oFfIqyMJKzi5yQIsTk9efdu+TLK66mKAcMFg
hfXb02/nrpQw01D1sBsJ9eUybLSMuXoDDeCZGhoFaQLuKGQ2BDQ6xvWqhMn2KxgTHcfnmkh5A1O7
MFDtWKUycXNHi3H/n+tq6jTtuDwJRpLe+E3KvwFFX85Kcmzl/oYE0L5HN0WzwJkwLNGSw0/KhsBy
DLsc4+p98LIEu4oGi91QJ4q0rpMEujOFPyJ4LTDbnSM38ktqpItDDRMZG7fUYjBHZ3ctbmpGIg6z
WLx50fPjOpeg6RQ9sgH9dcHeG3qrD60FN9dpPPEY9RQwyXWRnaZ5/qe86NAiv5vXEnDJRyKOP0ET
MYrL6uDBEGZlJoiqzvOO4OldG5rG1kIt9KlB4Rb3X7u7P2o7wfcCcaC3YnsIIJq6leLhcWJNYzH/
ChOqfbB+t93bqASVK84/e100nuMz0sG/BELJSNya5w94seVU2Rwo8hn6YlyUiqvkAX0TXwrQ5d9a
7OI7Yguw/vOhML/J29a8VvhyOGVN94/ckGCiJchcVhUp+yj27AzO3B4uMrTO0pMWF6Z/hT0iFr9v
yBshwTp0un8Y6Fx2uD/kjDXTb2Qv75hTpM+I+WXObWd8a2HqFScHEPclEQP2zmZjnvZSL1F3tNss
gbNF1PATFPXv4dFpx2HgMjyDu8J3zokZE2A4enNhfOZIRPgIWffesD7VD87U4sNq2izDNt3u9Rss
0ZzLJaMGimRjNJTTIP2dvsw7pi1e8juMkWlWzcHC+432nnMx54mGZ4qiq6TAj+Fes8gYy6pcT2lV
QDdxhOKr9pGFiGoz+PPeed5GtWLqZuxF7H2zoN/9GFt/maD0HquhvpkZkRZqgtJiDsQvrvlizQtx
bn1UNhZ98q4zFw3GACikkDrwKjv4QGEKDKUXzD9tQ6Io8kjBQ2KbZIUVi+jx/2geqdifR2ehvadb
uBbZAr41fnW+oUBmNQG6PpPwXs+Z9R+ZPgj+B4HAjJZGN3iT8wS0i4XBR3hc/uZgtfyEnZxLT7+S
aTTiiJNvPZjgeUqze3w0vxZ6VU/JI4Q+k9BPnW/rIpzrtjr3XzeQQwF2LkJbI1CJAnumONi4dZaQ
9emVl5aZ8MMk6sVfn0zUdkq8YFDupCcHB260z0gham26V041xQmlEgohRiJq5qhpgG+trcHLt28f
sbfVQhoni/K8n5ae3fKA43wYezxUQuW+DnrYiwu2xjzxrJ/VWvx4xpj1DNyveQk0e56bQOuRu81g
sTVliK3exOFoIF3sUAs2FBibMgJ6cOE47W2M9H3O/Q2BfLHyNz+FXwSmMVXRb4IGS/9wMhMuWF3a
j2HC88JZdNOsgfJzKPxV6nw9aYHFHQYbKQN9SNGpaNMMFx1rgKxFwL6NKNKZfa1kuQALNM7NtQEq
YRfj8c+Kj485czxGF/w2oYsnaIjT5cm/aQFg1ycuu/X2EoePizIIMA/AmbW19Jo/dPgeY8mZHGlm
3Oh/bwWgVI7JYh3RhSs3d9BwQzo4WHS/kEWBGildls03uE1RfdCM9NvJBTLYYsVUfW5lOrVv7FjZ
AjPO6WNeOA80KpadxbqsrAZJ94ZEMRh5DceMH68kijrsWAx/ys0s54rG5x5WsfPVbMPF7XUCoHaB
PreuGAWYFjlnWwyH13yeMDH7CEIBpHuNj1ANv7BlrDh/itsJEKZQXU6/U7k4HGHnhVhH/SH6V02B
isbIDvdaytoQSnH2qQhRXvTkSa4qUt5vpwgAQzXYOoWvfn+unQ6cBqkQP/cuoGjEgGjKBgbqk6ps
uBBByKY6QgjN181ZJjLpxT40FuZtlbTK4sM430yG6iLukYyJJ2V4Ro37Fj2kgr/fg4UWVgd9T0Nl
7UFlZayxk8voSuPVMojXDUu5QXIP3H414ZKf0cykyFCwycqgQSYZuwudPatZe7jcgVmHb/PXYqOl
PUVhiee51h2Cu9AI6Ejq0c8MkiMPpKiBdXRfYQcl7Lcwu0Ndw9jRvYm/dGxyf0q3a3jDNjapZ4CC
L/s5+9olUNN5RL/uFFQsQwrqylWVk4A4wlzZSDFA45Y3uAEuiXPEMHhrHiuCJ7rju1DyuoJzEUfz
mjURqubX3bK6Ms+0AEKmbf5HA5xzPrhF6L7TZki7pNngam4xFMXytsMlkMMSwE1Dz9IjCaip2oI8
rAOcI4Y/Tf2q2iKwQ++uVsog4lVhBxrFU4FSrbYBqgxSCi/YoaMV6S/gj9MONMBbSg10gNgeIegs
wYiPMInl9YTMKFkmGLp1N9lqctDXv7MG0CaxuT6vcPjY2KZ2ksRj+eQPAqaLvJQiG8FgjHl+O7i4
m9wsJ6a1weMGfzHYxYTmjgCsO+eotoLSTsvuRM6z/cGTqnsxQ2Ry1q+qMztRnckNe9lDxLw+l0p+
ry0wgjiEFX0PGo52KNa0yoGXNl9/9In1OYwseqY8gf1oHwahKwrcmUqU4wPbIo9yIRSEA3vHJgYw
Pmahgoe1B8JTgm/ZfUBL4SGo5EAY26bJkJDzoaAM6WEwclha0/TWWBvwkS8XPHHOtO7drRINmoiZ
wmiVNiwBc/42n0vjq9i5zZZ6UpTBEn/4QCWIEh7wppNjyMxj9x8vmEynveyV3SQZ7L6UIBOK0suB
0rHrYem3XgnBtVKp9zdal19JVmKC+t/r80vgSHXlBHuofJBaHKn4ipbmSaZX2U0WOodqWEmBuGcd
oAbmvKbwt3zL1sf5QjVvqJ9ozVSRDxRt8M8xP9ofUjSakVWpwFNx5/6yRcOro63yBkJXyWbxeQgj
kvlKIJFRetzDzRaNu8/Y+8waSz1mgVmJmAwKDtQJgQjmh4a0x6HQ97WDpDNTi5LBag9agjuHrUuB
ptjnaMMvgbnNoUkCxqlE4iMoo1gM7M3XaVBV1UT3aIkc4rMzGqfllMTiY/+3Dbr3S9749HmyO52S
azRZ21yGiEbEjb2NZreQUJhKubHffkBFHKN+ss/1J0D7euce7lXWPl80iSrEFfsHr5pssQozLTbz
kzI6xBOvUTb8S7+nkNLVcoyzitLD0V0rYoYTqXhgzQaEdbGpw1tyBbmA3lfKTrObVQ0VWZD/bEYH
mxKxEX1gpZsII57Ck6XgbXIJXirOqIj1JRfPY/KFE5mK74ubCNrZJCPZH/p0+bQRACWNWQWPn4gc
mj3X4qRR8otN+1iQDAb7cQKnHxgJ/qft+4vVO4irSb8fDlsetgPHXfMxmsUAXbiDjxhmKOmlZt45
SK8qyw4T1B2m5TpBoBSZ4NzeiGPalRlADcXa2jTBqarS25J9qpOdWqcNfJabNQRJ8NoJ9oRFTYLs
dvRtfC47/rRttdoxiU1XRivdgDq0PFkTZwJi0zt7+TrNl8/awV6njaexYJbW4pEsveuI452Zu7MM
KH4f6JQjgCWt9tHO7YtVoPoKW44Alrc82zz4jv+YR8kObYfGZalaF+GQGHoH/wjBJPOmvOKmNd9i
E+QgIepX2OOXagNmjCA9jH30HTWvZFssUdQjrSYLZU8xD6sx0MD3jBsVbUv57Re/P0CNU9kZoNfi
mNGUtWCUPn288NIOGZddEv60IeSHkCo695tTSFsMLSrF5hmB+qiHkPFsradi3GDbr5VL8kshMNRq
Y4tTk9jdUM4R4NKNRlOsay0ufOeYeCvS5hkg5+gp2kiCPqVjdaPZLlOqtnL5n3ONks0O3tMkxTme
pMHeqlwHmrZJEcySHjk+o0GKOaJwIdogfUVtC78BxV60bM9tEzFtwMpAA7UOHHEHm58XBhZpfVu6
l2Ops3sb86VC9TFAGAyBlz2mvqtx96nPBBCfEWisx9BUwoeOIcJ48qVhjKsjJOXwXtU2BYtnP6u0
cBd6FN4W3nWGHwK1DgUgCCOQPeYI9AiDeXunrfLg9JJBlGPG+HaKku0uBN71yY3OM57GSgit8d4T
vTvAJ7UbfPwUzd9kaEgSnH72Ax15J7X8AGelxew1GmKxD0XLUIvM/6h9ZwT7iLerIH1UnJopNnfp
gjM2Qi9hUUwntfg7Ultw6bBdNTA/KVKMX4hw/7QNZ9fdyZzvg+kRaiyb0C/mc6uH7L9f++DXwlds
pk53msnSv+c1bmZSl2mQw5c5hUKTcOV+PGRBFqkOj65Ox90E0uQ2exGhrtfPRoJam0rYH54/bJJB
bCq2JTENIhI7LQLJRuOjhXQCnFk4RxAG7maXZ3rbjeirqjsqK0vk8UX7EIiz1VA7Wdep8kTFhKBg
pipGbQrySBsRMaPyylcIoZJnhmRNLVapiHTYiEz5YbuIB2udO4PYFxvPFt47rM70EIRZ0+0SvD16
0caJ8vdv45q0mOBHFUtEllugtTh6rjZZpamOCjnMjzlWbatPq908Dpk3TcApVtrK7PGJV45UpG8J
Bj7qSyyK9X9XTHrVNr90i7BsaAmkVP667BKSoNzvarjJOPfFCskOQUfAN3brMwAsiBGG/rC0x6b0
LxUaJsXtm2ngENdW+X568PY2/UnMeezkOu3LfTMePU6Xp5pbDkCy3om6buaS3qtlfPL9ZFqioWmU
A2tuoW9R47fVO78Ucj8G1yWwH0FWZmiY2dw3TVKx0ht83jHIPLd98up19nP5yNqLAenE5P2shdA+
D4Bc5eEcvesgGw/z2X75oULrvCSnlScBu5NMXnC9lPAh+meLrDqlyQWoghNNgiL64UFR+qGJRA+A
EqAuuj7Aly6VJdtyayXEwsI1oHe8OZfOwMi2MQdwHKrxnHnKLsT1Ex+u0n9HQaZQR4bKDVe+JWDB
MjPXI1epG8Q3sV6O7l/kRyu6gFkd+Oc2HGMOQCGXUm6N72/G327gOdd21aURMNmWgUSw1cqz/JQW
uyJDvHFx/DFi7s7hhC3b3eQ37L1PG8V51ZBS1hp0dohW4H7wvwWKfhcZPNU9Adf/74djFgW0w9WT
vcH+ONJybTNexcRFTwb5PcmH5recLQxAMVAnrAjxVSrUHIyR3rj/YAyqdQOgdraCb0a4ZUE48Fi7
0uutxFLIk2sFdjc7TQUu2vAKKXfiO/6/aNKep40o6xH9zg5Farti5Qe/VeVTdVPtSvXUPk3LxN5n
6Wrx6JUj/mw1SmGx7ZSZSLOvILcdgfaHkzUx+M3T+dN0u12sc8A2dB3gmgJDDNJrE+KQmCxlOAo3
9YLI9x1TXjf9pm1vft8e1ettpeZHVlP1FvfxnKsn5OrXLwaLiH2QgTdg0jojYkfSxxNWeTk+GXqX
XvrdoxpS5aUryCZi6bCz/d5+ZtOw81qYxPFNK/eVRfb8400p+UbkrPueF5O9nj2Ou3YFl8TbfexX
0FO6MrCO/ak1qNapq7c1SQLi0RslO7GHavmOnOUs7VH+h3jEHMmDU9GRfc6dBm+JRAMBbDuNwCNZ
0zihbOUs+kSYof3S4abyz4q0R1n2cWHf15pzcg92VG1gBUyg+iGqgChA0Fod7Aq1BXn1PGcUQck1
oBRNZ6/UjdwUZd+NL5Ffr0T/KR5rXJBbe+70nHMj13Fs6uiEceZr+XeCE34Ht74mQv5Vli9oDPwx
ty7NDW0GW3GY+SsgLEEqQchHMIy0pbvennzcTkv4NEHAfr3G0wn1P7DPK9SXeR/IiCMa8pJG0hWy
CFsOoohXLd3drsYQ1l2ouN52/pYdmrFWngdjrxi0TtrUSmrLnoIIX9CuUWW8qX5FTOY4r+Jr4VUP
DlS/mS7ag2Oj+mm3mjvS+V4oKivVo1DzRQgfN3B9XZ26yZXKJBO1AOX4w2ZdeV1YxEXd4MPjCYYU
9uTuLTRaUaB9+RD20eciMrrrwqw/KashgEs44DeyvsfbmiRsswJoUbevR7aCgHuYVhmdN0s+TyLU
q4U9M6DZlIqzdyn8QDczvIWcXty5BZHUOr9UWlhG3D6bd8wJKkUAIJRz4gKwVXwwc+5b2Edcqgyn
ozbTEAerpCxeRJXW6MQw3k0sp2Kh8qIpTMOa0EelvcBA4TDvPbIm30dXXrCLvJ8fMedGij7pgbMF
+CtFGaZCpneDSg+5lGGNluQ+Fh/f5x9h6HUpXwVf3FTAtIUCfDJm/rytBN18eYc/oCjWClG9ZXqg
hYOEmybkD6RtQUA4MpzAYejR0hWCsX627eFUBFzmluchVRramwZn92U/weMTH59tZJXrcS4IYApQ
ECbXIc8vc2FkPZgYd0OG00wFsMu0l58ngiuSHGM6dCwzD7dAWoTpoPXMOnHAV4DV2hc8cyuqNzl0
trXiEQTXngzSz1Ygg9tI8AfFDiVei5IwiEyadRJ4TNNZ2w1G0IlDFw6x2DE2KISTmpiqiXj4CNq4
DFAru0GvByrJBMr9rRfKZk/ilKHVbVj8MhiwspPbHKRR3un1brMllgZ+Xt2tIkWCAeRzomACEXnS
msIxtiEDSH3pP1CklAkVCHhyDkoVtJHE1o/o2c4lBEg1qS6kzYIVaQ74zss36MWwHPrJW2tDnwsk
wZu2yoptQdkc5rZ1Cbdr/GTtSMpPwMpoK9/YLQ4pmQeWeVzoIZN4HxT39SeR2DmgER7ogUbJISgH
6/BGLtO/hsB8FW2ic371iPOtUXbO2YGO8Fl914IH/mt+dA9gUWlRcgpp0h8udqA/xdh9kaC0Lj2K
jyPMI1THF6XTH9MVy34YwdMBF0nnRIEDkp6q7SWjXmCRdt0O7fxRAvO+mEuag7S7lz+/D72AItGX
o1RwNas0WBqEwC2hE8crkRtVn8JkReaXsKX9SC3mm+e5ffoI3hUe2Mb8eP1fvAc7zWPVh6SZbRuQ
IrqNDzBbbS5w+OwLq+toy7x8maB7ro2TX70gGQrZIrISM9n6y1ynafD6AcHSDoXgiLCqAuwD0w9Q
OZmoA0KKUtrRT7raXekoYkjcxJgqzhUjX8LDsk2Z/p4Nx89X9JXgVV1SJQgZww0gVpHtab14/m23
UCpcV9W0iX8cI3PtRrp5DLXapUDYrqqSDxMsuP2r5XD8HCgHUDGx6BwDWy6+2XzRcD7khDgD/Pdt
UoYXhdohMmQUtyrqlC9SNae0/SGGg6CWCwyOY9I3ptjg7Ft/qjJFWvMG04hCRJfpDtzv6ba6eCFu
yKuEkUstEOH7k6xphtkKRroflOgDeo5tN1x47a52eqY1ix2Npj+CCqem16wJMBlAGSPIEYr8GGbW
w6FeYrhRBiwwaaIejRWJdpQNv+MjJ3YKW0dlEU629/SWDny+F3n+BSO+7YdpgbXWTYzqQpo509Dq
jmGC86vFVwEdiveQDP4qLTjqrss5xg/A7nB+0LzMOss98omuOkvvEe8laTJrk58pDaKVH8JsZbA9
LcEa7YMeanh1/+jt6hyoWZEelnEO013SHSjrS4kQYYqrWAEQpjceA/k8ZoI7jedXwJXw4V4KYkH9
fz7FuSF5CzkVGSu9ANDILsuG/OWs/827h7Z5OGDhWkJ74dBXtDpBfjbyolt04uqtWW2PSpPHVEjU
/EY2+9nsrPNhRpMaxfXZmqkYyBoD4TY49urOm4D1AIynNNGrFD2Bh+U1LigB0R5bRPFsUCtUzMla
8I61cQC33J97U1aWcPFcxU6hvJLzJccXlYrnZ9ssFtCND9G5K4ygkWUnaWrNImUFWMeG2nqkHmZb
WKHGpDkXiJfVCTUEoHF+YVpekCHovjhx+V6vyei23I7D/fmQN5vkAxkh7Vyzqo9aIf70TllZnmxC
6l98mSWFJL8fBymK5NxOgPYzcugw/HEL1WQJlJ1Bp/gevEvf8mntC1lFEesWVH6kniDvwXs7syUz
MOe6qREXPs/EU7ee6o7rtLl+ToR0B0PqThpxqYGW5CbbLKEFwQTiFKtX2XWNLxw1yJvbxOGwsA3u
2rWhDhs+ttibKEDN1HKt6/zVQXHR40ZrZUWjfokKphgyyQOCTVgjkX7udqlb8CTFcGWm2C19GoxM
PON7a620+KYkt6s0vuKHqZtMDmzDt8Mda17X4VPMWtE+XPjqF2BrJdw40LkIg3tZtXcZNUQora+6
jfESZksaoA5wKPpB5Kh8zULKBs7sU66TzIql9ft0u2doN8okl48F+Zkx4LfCkuYvHvGJDKxSE+Cy
hE3m9z3C4au5uIaOT1XT9EvmrI1UgZptvUWtGhZNUb+6H7EHo1v5X5PtgqcikeUpx95LfDdj+lUO
+Y37lUG/7HtDYDn8iXba8p75XBsohSNUAdUM/4dNC9LEMQvIpZy8wfWA4ULQp+QGLSE/+AO/8Hs1
Md95iINbLW94TgOjRsanzUHTWh5ydeDdJ2Ytj8vpdIoZOyNYQNurC85JrunRwdiBk+yesmunom93
OBm6Ooxhf5nBC79VlyFUoZPTMPGYCK7Czv0J4TcI4u5jfgHYaKbj5qPPiAmDowhc65DZmSRqLst9
9Fv8xb8rzuZAbF464QE4wAp09nHLeilnZk2hOadKGML4ixvhfofocxA/e8alyn+LN0zxmfUPS9wW
/joi5GXBhTcODJCHAbEpt5ae9k36frLBByX7sWYTTr8qdU3akl7yGzCWHgtX/8q2mcuRWj+Hu2FT
GvewyaVlF6fSOc6Jh/ZoglxtVXcIpy+4trGGPnY2suS8t6LBYwAaNnV7p2G+56ZaVwLs9ATiTYHH
cVdSJECxMWKozXeKtcQK90Y6yQimLpNWFoLrPQ+cux7I3anHdvcS1Dc+FX6SOPOldHMYzwsx9vmq
BhOlqE/ot4aDF6VoF+YGrzTXJxMWH3rPElt5wcPJFiQHDFeRM2OlrYRHoA6iatkK2uUJ7MgT2RfU
RuhxDnThtt6aDD2DVrv+pHQY70Z6tB10ZY7rswhfxIcsbRQmPDBqSZHflLkAcmBw6aAImLqYyiDb
/0ty9SxQKf2a4G9IBrg++EUI743kfWYw/4tXmHb0WgyBeO4ObVlTCE+rjqOEzH3rToEXRHCuIZIl
3zrFFR71Bl94toXigKnt4CvKx6htp49/euM41X7X8OM9VCelqpID2YWeWrpdNnR0JKyAnlc1tLAD
z+k151LdB4IE/3+Y4xHOlQfYETW0NIealaMA3S8/N1ifky5w+cJ/xonhibE9sv07XF4WyekD3TF3
243/thzciXEaMhgbwlbqt31Ypqut/LTBaQ8WvmQw3af+muEHERops4GzAF7Xv5R+0GuUPsVRgzzD
ilVh5vfHatEmndsoLmGWVSV0z8dCIMpdVxcQydEb85sZsgXpNsCi1XjewG0u+M3cVGun1Ha0G9nN
1hOhU/kvd0yVSa/04HjPPZQb+g11wBb9WJSYredQj28N4XcskWIj5nPp/bC115e9AkM7e4P067TQ
33qHR4UPKmrQ7zEFF0IQWaXLHATEKjU4PQe9vEe7VTHnsgKogRZ4u/GlVlvguJ+E0gutci9Ii3DC
5wcAhZTkcAMdUf8gDypTSif44XX3APnvgDXORiLlACmbSuiuXcRJT2+dZwVZZHB7Dm9mvS0Ev6ts
HlnJA8tsLXRRS9YkYSGnzhdf4W7iKMmPN4eplHS6bPqGAmcJEoi/xr8K/RKiE4t/dprl+Q16QAT+
B/rcyVedS4FdV4yqtY6A/1/VTkiyiL/XHHAfm+eZxe/TvbEYYf7/bgCbSJpehBTYHvo+c6UbDxyD
ppg4fqT86fDxpVwPOpIQfa6QrT9S+QwSC1zx6m76aHIzyuF4kGLdSunYgcfCFLv3etjRTnzT+eh3
owe9UTm1l7vBnELISwmL4EL0XRXfTK52kZjb7raZN6kCXhYNKzYB+4GG0CVqI7DXZMiDilV48BcE
aK7hqvUULPBotYCi7qdSZFVGpkDu2kVD36Q9NBZpBuaUlxjobUbY3J30GNiagZbn6NFDRrgb5GXM
0PFXEsAViilNd0/LhF9KVa39DOjFq5eVFDL8Lw5At7SMoT/LSmlco6ZsweTZncQEXdyXwOBi0cl1
uzey5qcJPtUI0tgqvPANZxmNulRNRcbSbW49LD21Fs61qJcRjuQdhuKJsy80N4qDDyG+E2Phqv65
FLwXKNyco15dppCewpnzLzhQuTWeFlXJQZ8o/iseLce95ARh83DswS2BVd2MwtwUqJfs7Qc9kjb3
Qkrf2/yUnu73aAZ8UvlCRaH6WT8jsDm3SEBA+4+KlyQu0jEEKCSnLL2KLkTbCbQL7+pDaSWqA+sk
OwJ7mnFUGSL6vsMj+GEQu86FeaCoXselOu62bA7+vuguiPetsskxrJnJlZ20QpZoLwTb8BbWF82r
PEMETNMGRLKM5LJzk3vJeMLmEh0/vVmiENrn6m9EoZ7ED8LFW0Z6x1m4YSA6q3vbCFrwMzttQgO5
SHuPYMbaJZMIK/9wUEosyHhKiKurQccT5WZy19O3V9/rKPp1DFiImSTv9w360h+8EyFZa4+ww8iY
Ao+DEj7a2+SlBCDDuJBXyqzPn0GGf64o0Rg/JKWutmyLWEpB/on5dZltwHPFsJuSYADdNqTOKINC
EMtO6z44e9bJDDz380LF7Wi2lXC0EIXY/F3T1ETUMN22f1lD//wyf4SB35wZKQdq0TbHohdvnOi3
iS+OFai5CRX9g6dkkSOwPy85kdQRLv/4YEwXNMfQDLV+ktJGgZ3/4Ca0VMg3A5j130B7MVY0uNd3
w1cCLbeqhRALpMi3/Iae6HItxwRdwdM8dc9Ssdt1Q1S94L8ejMaZilhpLTRA8fQAuA1SUMpS69Au
mj5AkMboSUUlEENvkVLlGh9ccfVsnp3nNmqHHcOo1F8DcocCmQDeMaz2I7BWOgFFUFD2WZs51mMl
hzUs16e/KLoP1KVTV9hNaSmL0W9g/fMOsnQu5/VMv2R2ufQpHv2SVYgJ2BT5cLuNCZEFA3JO4+3T
D0ZDmPvQOImFMKGD+75ERSM1EQa3geLjm3bHDlDQi8cfYzb05GG8yZPOUlyxyLwkITMiq5gfTIGz
gk0aUTnMYWUtJoatEx6Pq1wWloKtgJeOfyJe8DmCjL5P6x99C+I6BDAVxeIVCVIcmoy0/oo20Apa
xV0E9wQ38NnQRAAW74Hx3hzp3z02330Z1B+VSxp23/2rH85aoFaZP9nt0Eu7D/C+dPAnK4oK5b8V
3n+wOazY0ktIbsyz2Kb2fcbMHPBXXWBTKPEXVBCUr8PrLkWql5Lbuinmz8i/sJYWlYxSCl+P8/8R
krUDJc+s6k5zQkhtR0uxEZgQM4FZ97u5QE358Got/PJ8Y0WKHDvVczjzlVz7dhC17fGI83GZNFQq
vN9l9TlahHHtsOCBrijLTsSh4kBmnkSW6pm+P07DGrZIPn2UBvSrjBXAdd8AFpN9ejRBKYqUBsGn
YPajp/+6zQWm5YaChoRIt86+NOVIWOEdlNyagSQsCct6/mg0I0FoyrPukCCTviWZ1nSdWINBbVJH
/SaHp/zofSBFko99Bmu1jCDftEuuNdkQ80vBK3vHZGs6SzkgFi/9uvU0UVXHlWPUaZCV2PzaZ4fa
5PTnjxeJAxMYNDSdRTta3ogJbThxpplqKcTXpQQMIHCuhz8SkGoMzeLW0/D1tfxAUeC2Cb2F1UGW
ZNghGOBwT+lCg2LRdJ4Ct+YdoHFQsc02XMj7uvZnfW/9a3bG9tXmSnr4p08F/f4R3OdOIvZUUZH3
HKi3TMYugPO8hpFrZzqAorhUs0UY9eGztpSd+E2Y6xcAWPSQeL93AaIBcV4j/MJ8Sa3rGYcFHuZO
jgK1fPOOEWT2C4C50vSwqiye4jiEbhFSDR1OJegMG8gAQZhNhCZY1I8UTTLkKSEaPxpSN42Yaa8x
RV0XLHhlP8mXm25StHbNU96rEcTHhCSPuj8mMnY/ZxmMWEhMkei8kBV81QaJ5iJwHv/ZSfPAzRuz
43gpRsl/Icasd+efZTcsAnvF1fYFURyDTvNhImhe+vFqUhZ6pW6PN7L7wO6PmsMGvU4tgODO88Bo
nauEfgioEZR0MIri6Ek3reQm9oRj/6XNKe8MhjahJ3ndzcjrgRtyKRt8dwBlw5xKpK6yXifDC1un
PHPk/wjBN6avUo41Eufl0qYDHHQo2rsyXFg9cOCngU0PBO/+9ezHgB1B677W8pS65moRfSkSiyFu
fiTJru+DKaj3+WQTAXiUcAYHlzCrXhwft9yF20k772zvpzESzT1+K0y75FfELZuE1T315Xa0QQEK
v3eKgGeeQK37h4JyNXQdJ0Er+GO5DS4yJsyaipJ73/C6uaosaBM5Vnr/JQqsmiiyNNniYyyt0EAb
tWIWRtqgCMN+khyai/1tHcfEMAwEm8MnZ5NlvAs/MEbpKK8B2IT45ttyrFM44wsGVhxdaerQaRJl
NQJGkNZmfferEKlYbTk5JXFwcmizRSP2wNjtqOUGzDLy8EF1BRQT/RPLnVUx71/MpWzs3nb8ZyPW
PbUDQKH4pKDB1BYe1jJlfy56gv3YjbyNXhPkmMZglUwZxaC/leCtF/wHFupKCXZ3vNqGxt7vg4Le
xFGtL3BLVFcta5A1lEaYLSl21iCoodaemKpaNsLTZhDuRYmlcS+FDWIqybEJKg5W8XnspQhzmPlO
hxZz3qR4JYIaCA/1e3eMBtb2Sdt0oImzuwZw9gpEOGDhp8Ncx9LztHcOip6bsbAnP7EcQioJHEwZ
VT8gkbsvBegoN7FCpmXWNJmvTrmCQl8B1xgyZ1yu5A+nxzqKOa+3jur6e/pVJV8/nt/nZmB+ozfQ
0HxDSqCykRwf6tK0QQ5gdAcK5UIpuWhKWDiJI4LkUoWN7YFl52NqL0aqo7lpzdePRZOAM+nSkCcH
8fXR0vD0vvMHBAvNMXi4fG0ckzK+6qb0iU/ktHNsDkux9XD9MS2iOWCha0ESRqFkKvQj64EU7kfa
0fw50tGUkrBnP9ktKgZyV6ywBqY7V1XxEVsbvLWSlLiUvIqcCX/YG33fdEKZ/s50J24BiPHiCDV4
Zgd9OSwtFXcwJIKSg3Ds8Z7yTsvHK2JNDyeoIfl24/fbGJsCGfuCCJvJ7tMCDadwZm3O+XaB8MuA
q4Mr5bh9CUGbLibhlXGX5q/k6+GT3inTh/YgeVRm192Heq4eybCqrgPoByPH81khJKm0LXVVWD8V
WIhHU2zERHbC6l9ye7+PQMX9AoRQgC0dY1rquDpi9lPeU7PtxHNcbdulVl2pg6MX9xmnzuK0Pd2x
/6k1draeYpCoHQgZkUZlbWqznJI+RkwMnEUk2tVSQDvvy7xNhak/eOpIvliiclOR5vZNQirXp8+S
kLZZ65I1w8e7Wc6vzRg5lyZyA7LtqmG/ipIMEIhKC0kMj+AFRhoUnRPHf5PHKjBHFqmLNvMRADDZ
ukdiODDG0l6go33251ifF7Ee5ugnxlNmveLzL542RRS8Ez3ixYbfJxqmqnonpj2Vh03ZokDGrsUI
PNbMEuwZ0EEsru3XpTEQSIUz9ejpW5lYv0ZG74cfjY/kc57mszDf8pGjUhH6fkKExww9wgSbge42
g0ByvM7yVlvJRFowisrG8VartCRCDkwKmxnSXI3i404luAe28jRDI/YedX1HlGzne2mUGEhlSxZj
vUk+TyaaCLBUxQph8UZrO+S1gnBCvNl4pthljSDDF0YHbYUyBjS69ENYPJsrGmhUMLR3/pUpdCF5
b8HbyvwSPYSmaORp7lATfkbWZIBiPzm9xQz5312jqVGXZm9wazNC+AKrMCSShAkDZSYZvcTYlIFD
S4ymEIOWw1tyEwqdw+cbXlAVgQ7NxFhEzYLQT7TBWy19059mtjKWszPjHJE7xEvUOszNYJ5ikDg9
C6BYpZzwQLX2TsqXmq+1+eRp/YKjIPYJA7zD4jNKY0UIAzPIRqh/9zgl+zfEU1+9iEqYPXOONFrE
WRDa3JXdhQ7Yl4TdOgNLx7MPrANO4LAAcm2ruAYiv+CL5K6acS9pSfiM8NzQ70LyfvgEoVmWkdnb
Ws+WGzM0uVPVcs8MkkSdmaAJHQuYtEOTzUxNQ/eAkGQOknf4xXNndGWNat/l+QCXYFnRFJPe/zUA
Ei3YRW0WIizFvk6hCwQ6PKy4DAW7KzU5jgv7MMG4VvF6duOh6cnspS+dxhlgZKJe+69Xv1jQyikY
5Qgn3mLs983GCAs5YdOMyRP5rua3FLNLWcbuUFP48HUrM0B2pt8DAhqTCQrOdyRibzHqCKve+R86
hnaxGLUBSOh5BaLiQkyemw6Y7Qvx967c3sShxQm9PvEryfYR/sWITIjjTdkYC0HTNF1w+Dfv9EaV
MGduV0xkrAlRHPM6gJS83nNW9jf14jwebJoDplfslqzOIW1xUeEcdEGJDtjTdEeCdTay7pd+2Is5
3L1cmXhG53FOLKSJdWuJp3Ci+fxjjMwW6AdkvgY8+51X7nfHQNT3fM6OjlpntOtGCTwLeQU4Nq98
H03p+05X53PNtUg5HN7CPFHBhp7lCyBpyelmlVLoiu2UITXZ9Un/XBl+8YkWAvOv0STpy0HSic3g
6EmLznMgqATxvtku5M+2wZ22hnx4Tr3/knJwEwwF9LyDiWFSwRySAeB9FwS9GF3nhJB/ixDJ/WOr
8NVBjx6vi6KPJyEZgH2Lm3QHm/RE02J+XN4cswDTqhff0MSDHdXivETRFqYRM8gBFfcvsYlrf0Yq
ooN+xRqdWSeNlX4kACOwfqWL3jI27RIw6OCOUpQmvAVGj/ZswESoGl+BInm5CdOc3B6sETC6oUxm
tl8lV8SzELeatsUhdakkKYvntVZWvIekyYGBUahatra/ess7xYGqNEqR1LAGv3QMxrmyS4a1pJDc
550DqgyjuxBzrkNuHevFNUp6KxBL7UncEnvpKOPdUPvvbPQNwE/r0cXxx0m2bIh5XnS1YgN/SDtF
5dMw1K5BzFQCN7xITHgfMp0Mqt6STW7iq/wVF6od/5a8yw9jm9y7GYaaudklkvrfDh1FojZjStqY
hG5RsAfbYup4DFQgfxHth9lKy0XsxfpOIxtCcf63+vnlqaEtOtOnNt6GOwc07/eRfgasjroOJD6v
T+kUoLKxTEwLPoDOpuA4uP46MXFEDqqI1Z5D4FwQWPnPuR9ewE+zNT+3/uacw9DrGSOWejiAnji3
dayLNT2Ufk+DCBmeQCg8A1Sbg2C6cXaHa5J6ub8lX55/ei/dqyDqE7Ot51BepFl4Y+VZLGOAfX5Y
mjGwwNUj5oQXyFqJ/4A30YDtxtII5Q6Qlj/LYsLOFYR2vkNn46j5Ghfja6iZLNi7Cw4CRRLZ+Ru+
J0MMEK/oZEVUCqnN8PdYpNS4+iICHRJWOlAjxNCriHKZXy4iCI4f4G8b9wFkk0dQXS99wtRrVceQ
Sxqeh6/dW9gbUsUySwJc6lO6Wt5s4dvE1209cD1rIB9Yb8SPGwCHjaPp7ko3uakci8i8Vv9p769w
7Hfu7JfSGloXCze1ksi8trJWI7A+jytWvjj+YIwIQRy3maai7nLcq6CD2s9KwrjQCrfrn8Bro6KQ
VJiKTQzwWrLad7PsmX6ObLQP1l6uggMUQ260k22J/+SRuC4C5YO41orMDIbsuFtWhHNmB+XzAscT
WqaGUAQzNz6loRBx0mFvqrHYmCbqaBLsOnq3+294cZ+tvLQmg9TXX0Wl9aeb/9kEznDKIlSpLBqq
P3p4YbGcZo0PR2X2KkEQc/OAtNp0++it+YTavD1G2zm1sAgDKZndxBmzj8J/KYN9RCPeHI3EqpLU
3dPGDw2GOs2TyBaSdXxyJ/qgMTInOouBPob5Ua6Q2xgJ5I8YESqS9aNsuDUb/ESz3Xp4hwnWvwZ5
MX83L9VmNmR1YLbmukg1oWlaVnui+GE+s/Zg81pmYH/nq7M2Vf5epAK8+qh93l5+fhCtPaS33wqu
isG++wIt+aD+I2waj0S1fZzzrz5p2ATl7N7FwAW10kCBckVjh0nqoDcy7K3OlMQZYqxOd6xnvgvd
b/xgDcTwwUt/MYAeoYdy9/EIb3mV8/9ZMn4+F1RqKpuHq5MuBFgxnjSjc16UY7cr+sL7PEmSFFdQ
vtR36rZ2+BK1wZ+l6iBr40oUQ417WUxxPm6eT+8m7U3cZQA/Rd0gdCKIvGfffDVvK9VxPxEmp7lP
jvsoU304xMoPHEAZzi9iu4j9mA6/m+dPjDBMQ6s/m6AqYa8DgXQ6/m3n8Ad+Hr4vK6bHkVEYF9z3
9q+sCkbYwNlQ1H4ehtVoXBXYXjFskkCEmAxIuoOHRIeWmoOEZ63S4i04mKBeE4j6pmwQ2A4vdQIq
Vuav7y4M+Qhwovy4Htg31XL+EBAH0/PybtWeZG9p+4i/hXaA96lNmoVJRtq6OCHF6VoV+zDCEu1H
tWjTtZmpMrriNsviPFyebVLfkd+A1QlvoswB4swyhEqpxHoM9Y4OtVa8j6T4up+Xk4PDyrFLCwRi
LRqPQmidWuXvDuAfVvvAyPZn6JklPJD4Iz5jgLnP88H31dwI8q3jwemma2so1N0O4CwrobkuUnlP
doYmbuZIo62AX++Dh9UOlSyNRCZvDnViShxXTk8wj8dRrwzN3vp95Pkpbp8Pm5e7Mi1IpJmm60NL
6+CnYQrWB7b9SV8FblxPWLV4n7/qTRp72xIhIJ7R9er8LWa7yJz8qdgaMx3x/hOMgqZklUdhGJ1t
RCIdcumcTiKbSnJzQ9kJpuH8xW6WXb8hJlxL1f+tozGDBohNaG92F7QRrZcXOH7NCYKjFgd5lBhP
SkEBiVJlbvn+W9svTzOa3EGCoKaTXjd5HSNhHME0hC5sFIUTUmEXptp5tXNrzAFPuRPqeM9kepsp
SolB27FJmtmT6+i8Rs27U0krrwHHwPn4vFDrGrt+nV8QhyrO8R5emwpOSDhRgQMICmEFyVOg8c+Q
PVjmTy4sEk8mpjBxySyP+BBzRzopnw4feDfT6klT7NJR7QBc8go2CRw8tK/S+C+sEsOQBT3CGOnN
EoXZ69rZnd8hMBF0H0qg39Wf6p2xFuAlzMJalk8+wkUCI1vxapcmWAtoo+/wA9l3k/1QpSJ9kFJq
g7Dc0th0sdHgGFAbdrbxfK31u5f8r1Ahq6oocs0Z7LEutN3FfErZzxzU3FjzqbTudKc0zM0leGH/
dPIXPXZQ8OjExr+RnBnlFMmyiKznEZ71anMt4t4ISjBLQyBjkLHCCj5mA3foVH6IRPgv/qksLKhD
NKogcKWsnKYwhkwveHGihlyXYS+v6syymg/yDv91krIADQfMAQIiUzbcRahUFmck3AAEJlVzu5N9
TNCfXTggfgVlKywoUkzeKf6YjGGYTwxu8t/hfkuuEjQW3wZuUFkpm3d2uxiW4m+BS7RUl3HY5XZP
O1c/deIMQ8hE+Toen5Gkd4IDK7dzuf0jrLDAvsTzKB6VAR6wQZkJ3JEqKWROyWZ6VFdzrFzD1Znh
4ysP728waqL6O17aMTS3EXpebr77l9hx9mwz7RzPBwkj3wCR/hKGJwnaOzxfl4FyjFQTQfgGG+bt
Dw86Z3jO96sYIHuwoe/yCySJv+VUe7dfxjZWnUrW1GEbNjXUHtas9qAV+QaS5V93ronoNh/Jlvou
Bh59O6dAQ0me/KcGmbTMc9kJXdeY4ZEYDWMLm89ZqsLlmv8utbamZfBfAyEEJKWJMe7smXWyYM7o
RNl4tmRO0wrQ+1+e5MtgTq52Q+N5iKXCgKlAmicFQHaFB1CLh15KEagH30+zqT9NNBo48f7cIzAH
pkuAocvbYb++/8x6I0DVGo1CLGphf4yqdFePm0KoJGh7Hqtzg8BRYawmXcSrTdEwaJg7H6IPJjSL
5ErzSelp3a2hvnCXE8zBaFTjurNNvBUCF5ykJaqu/FWJ/LNzrlYy79oBtua4fGSynmtj3x/UN7mQ
jTWcXdin9zRZSEiWbu2zwYCIAQnNLMn+bztKlccqMNaTVav0rqHduDDV05iw6iraOSn94VVTlWVz
6N6iPNamjalm2t35EDWZdpKn4QBoT7/83Abt7aKHZXlOuXmya541b1wAkymt7nsNWVAOm1WW/N3T
V21wUJyQaRvHFKcTWAnTSPqGMDvGEmIIOuJqq95uza9UBC1oza8sX68lNdFa2QI9K+8fBdT4m6mi
bW1Wejnfc9pXyfRXHgyOBMvu7YF5OILG1OUVuwvKgbs7dwgF57F81iji2ttUFgNySj/lBtMr64Fu
7ps+013t/UzY1hsZO/geXmS6FdF9HUE3ZDM8euOjIuea2vJQPuD4Spdwn/GeyY/sg0RIrC9ouMJm
ENbAhq9WDNN5IYdGUHkIVGgEqInap41KWwcmUwpNtlXO9f3aoXCt4XDqDmqfpnHIKCJlRnCGsKSF
AdAr+bJbuorrKOW0dEZsPRvNZcXwpo/G7G8Zw5zjREi1gAJ0f/Gqci0+tkWH1GKL2c3xpOx7fWPx
8Yi5PfA+/O898Srldg9zKNaKNcLRdcnWSD21MvUKb/N6BJgbuHkSFWMDa+GRmUerM8+MnDXzplKz
Ll4kysi7A4fkIgh8KARZiAJAFin/gvuv3/qVAoSo0J3BzSNjVeoWSSp1TcFwVQsvwAYymoPMFKeg
OAUYSQu83CqTfv1NO/yQ5es51yYxJMPFojezHa9wbeT8a7pCaGkF/cds7oB0kteP85q44bAqj1Je
rrFKY8PFdZH2h+0NvLJCq7Sb8cECtMWFv3fwOj4fXPPkrCrfVaJa4FmmVLk5c/Sp2hv5SwaxsiGY
VOQzexp6DEhUh6vh6rNwgc/x/Ls5juX4TeiCGkvf5VrQ7ZRciiX9DsXiozJYRaPYyBr/S78xp3/3
3XXuZm51wbz0xJunlm46CI4T2/Z0Og7P4nKaMKHWIZ7EEKZqu3+pfmzELa29PaTetmgncaQhL0DK
Hxfb+NpDQPGifTLE42eGs3H5UrNTsrYL5HlyRWpAxyYBcAkvyyKsKPz8QaMD6NSSu39YHkH63/JR
MCFGpe0TueoLA3lLjR1Z3yVIpsLqnx87pF3ic19RVesTtu5X5XDQmSArVqGS39bNWwavaDJP/QXK
Zy03Kus3eQfPlnZWc2MZnHto/25YnmuPKP5qCKvELfW0CfTIxLBMH1JH7fJ++jLCjKxZI0XXPGbA
4Wc8HFY+HH81iTfgtAyLpRwSFiZy0J+Z/8PyN0gEorNVu93xFwkIr9AJ3FSX4rWI/pVfq5ObE4sx
3HTXUz7ZdnkrOMgSb6AVjZSNDV7NrSJN4L2UpAQzyvg1pqUGQ9sK4fcFa1s22MiVaunzKi/vyjdq
doaiU3p8+1bdTk8LZ7ANV+qn/trMJ5la1OXqStCf7LHSqUxEkLLFXXDR9+ydIMD8eBEtROk2bHGd
fWJ9kaUh4VpKlz/wrOY11ZguuAs0IawqF0bRYQLLdWPyQU8ynytpNsANft8ezmWX0Yb7ALPjJC9N
WwKVk0kRrGi3cjO1pFptAgFfNWTE8VXK4RNMSHs879ylCzExvODUXKx2qSdJWvAgdYwselgSmZuI
9EDQTVApFIFU0zClg+Zai7IRjYfrUr85752sF1pej0CYFQvVKLS9muxqNXO2DC7UFPJZtbKdm52L
h2uFhoxiSCgdWcZ2utc9v6QePBsISg7gTvW9M2nz4y5iBCWELu8azqFv1Qt9hZOLHpyJTM9L1mIn
J4YL1GFjcafx4ARfwUrsL+SQpKYiIsWX0wnN/wMOPoVuIUBkpidWJyA3JbYAsM9n8oWe55yA5G2i
de6CXl/0jkCSbdhlawyrAUdpz+Fw+tGFQJhiGqNdenBq14UDLYLC4N2owPne50IFEftYz22qXbaG
cYE17ziHdbLjFz5K/5047RAl27X3QqZgKI8ie0aEZfmSmRZpQ/sYHBbpR7/vCZ5er88aAWrYKlAt
AMZGu7YYk/I1ZseDvgQBWIekUhhlEtJ0qbXks4w0qJsql8C2nLsl9616lY9fqWayueMBDwSGrWwL
AgX+0FWA1DxmM5t6/ylUjncRL3TdEDnE1maHJJcdQ9IuGDfh4XVvC3iNrGunQAg6n757mM3K0VIN
plb9t+1AELbhgxB1siWzX99K7Y8/z/6pqs6h3oFxe86lsZdAn4T6LX5lpJ/lvzNJ6AQC8/LFFd63
auVzqVIyn3XG372m/oynhXh4XgVU2UAvTLsI0ab4l5QDnlSueohOS7y6R/MZZFm0KUWPJgU6xeuy
AifRWHY1RdQcvjq9qYSJlIrsk+l54FwhaMEZ9wjS7FMlXrP7d5JOVBK1auXEwyN9Hxkfapt6E+ZG
l6xOcArh4agiEaSu0O/okgReLou0Z81Y3Llg7rL8jRAun8pxBums7O/TJUe/3rWQPvWl5/up+hYK
hlBpB0kjb4ocREVOSQfU5napLO/uugTnYJCLKpvFgQDJnowTmegjcrm97kwpAnL5NbixmEd0v9cG
QRQz0KdWIg8GC+Sx9J1KC/a4oeWETrj3mqcqNA8OCPgUWtqV+cptt6GAlb/dB/64JT4jeht6qaAd
5w4qysC8jg05qC/A7ut2CSac+4z3SirlcM+b1Ng7aMMdHnd+5F8EKVUm/5J1WbQRxvyWxDN6Jmw+
KVc4XL4P2cvxnqy/kPBvg2gtR6EScW/hA/TTS1vnt7Np0tmMsodY7FqirrXmSKmtWsPwbNKq9VWP
QMMa6Uq/FgfyDX7WfxEvxsd7QSKWtgR0Wy1ZLKcICDwymbTlJcqQuNzhwNPe1Kwkp3NU8qee/mVc
Dx/XSZAURp9DOlhRc+FOzGWPR6dDN2YDif8vcuqGGBLVw70WZ28igO6yYn8Vzd6lnAS0hTSmnq5q
ZDKGmFevsYauhLdLNW/r7N4hrU8gNHyhSVjDneSxXnM5ECQXqE2CrGfAyt/up6w/mkl2G5So/t2H
J4dxDFZLOzTmvXj+wy6ETJCZ8ZZZlArlVVLZybgfDfvRU52zlyygOUE/ep9w+g4lcxAjCfTEIQM8
+kredzBuAHEelyajdG14lDejCeRTewW1mdPAwJjtMwZicGWc8e9qUZFvWeCVQRzrnjGuThCdFNLP
Y/XUTz/fBotoWWW0CIRb88zebyUPnHp/KAfosYc72zorG6j/O5BrgnJUFgIrZrTq9W790KGC4MXz
xY7o8C79aKVWBk1JufRr5PDczNK0jUWyknVm+GtGudBNPvGlcHfVRObzD72V++l3BRCl0DipM7Fj
xRU5w5W9m9WkiPrxgQQMBHYxQU/ClRAtvBVNZTfYSgDzlYChNcuN4QB8PlstOAVp8WH2aJdt538b
Zj9xgbyEdVcMyzMojPSQL33i4ebYSZw4/LjLzclK+nHHUFNg5g77fZ+zR6zEv30PeHLPP9xPZo/O
dCjbiSPmdA+C6R/AfHkZM0TSaPuOXL6vdw+CCIdrF/N/Jdg9ciTSz11FrVSxA7Fx8/rrLWw2nkBj
C6VlPnXuRjiAdBTpIZfhwFwRZbALScVfWOWLsBLKo7vPT73U7uNUqxlIWZORYE4krIVdqjh8AhOb
NfpDQryy96Q+q8fo4PnfnuRX3fW/Unb4r0t1LomQMEi9DI22Ffr7OmfXDQbTPc9SfWCIT+zo0Fjn
1nyuD3BDVjcaHKlm7I08YQVo3rBJ+cPsRgE0eucOHESPhvmv7RLoUanvDBWFRZxnXxy+jpde2g4a
MzT+Z/Pxkq0Naqwg7IoHFfJB3vjJ/Ot0KIQydT5AS38NWig2Cypquo6TNDa3eXpNc8wXQZJkLShG
cdRValdVk3ub3nVBKMa2Y691YC7nmLXQi6vC4WI8idHXr0L8M7FtUPMwWSDkbaGNEAFoiFyw8AXc
MUmUE29T0RCph1lF52hF67OmUqxGr+ykMB5IQh6ygkYSQXHdDYbLAVCdG9nd3wqlWi2APY/NbPeW
eB/hBfkPydMOBuV5c88eKVEyXamM6D1YwKCczY6OPhVRtQHU4GWD24CSGpIWVdlHpOd9BMSts4fp
EHyvKLSITHNOlWx4sqwVsgwy4btO7lqxS/sKrGceMmrWZ3Y76RhE7/2E7L9Ro1FNSLIVSXnq0ihh
v6q4wwPzGx6IMyU87gUKfaFCx1xX+kbVbYjgty8JmmSWgVRnqmZ2UdTxvuebrYkvvE9po1SnSHst
/zmBooU6dH0SD3WWpkl7EY0deelF6pUga8rs1A1K0nNQ2kLuh9MIWcQkMt9zK2MkfdS3cjB6a979
6jJQb7gn91s19P/mUVWXchor+ikk0x9FIAVkYqVg78Twci+1sPoyAW5SYpFyBlrmTy9XmbnfVtuu
oNo6ZaYw2aYafiAJqS93wVObs4C+uClrL0ZatjwcWEMSN1FYvRrXTLBh0WqIrJuZMWi0Og2HNZ3M
6pGQD1vhB12JxNszIi6RW3B1wKa1NkSpAhoVJGFYOCysxvXMg4wFxYvepkT+KwbypiO4fErzGk+I
MSqyZVSX3aKKSuoIoR8i+MirdMSV35g9gpt86I2RtBwwzBmdnRL6ULj+7TmfJf81f1FSm6MII3oO
zsX5eokbutcijSplVZN/QFeFBy2IURlgDrXwoRy88Dxhrw2CZ7tR43prCnO74PYBVs2LPrhlJiMu
tfYQv1oiK63ysyJ9j8qSmxQCLwYV8jqXTAH0wzrVp/EczEFdQ9WfbX9UB1mw97UzSz3z94oup3FI
sgsB3AGdesN6r/geQ2He+RgwrZ5l3ApGlJ/aQeDioWRgX4gSOVKFXA+vU2pNU+BKQNkCxctDcVlx
dPrw0IULAVZocTx/C4GIlOcfX1TaPkk9vIykPDZkjAKmZJpudeZELgHZF3UyMV4qtyOn3St3eUkx
wVndHf5qqT312D6++eepulxeZ73/epilCA/+XHPnI1MamEfL7GaSuCsoH6lIe2MrcVSYvffF330x
/N+Ivt9LZVfwDSYugH7/0f9z/UtJ5mrHQAJU3Tdp+9bHgwb4VZeHu5m5vdDdU4REEAntz5VebOlj
7ckYifZtnEeWe3m3yJhQTW2tQ9SyyIXzui+QfsgXo3Zca+9cTto5Dyswqqdb2yx3unz90AnRYBkm
6efRybu+0BOgdFSt1ZlZWGUki0/d6EUhMWDftyWzSOaVADDhr8M7MBasmfIfGl7Alzj3OrLg2do1
ZLLikqUVg29dH5I2aSIY821WGXToZFQs15I7a5RRfftXtbyDAbi4Az5WBpEy1uX+qAfx/mHGekan
agnabcC+P/Tk9/W340951mlRBkZ5CSZpB2QF9htuHXRkxiFOb0kOiUoaxqk9C+jyAhHJsPfiymgg
ESv/mqqOE1fvm3BwS37nbawFvRsDiu10gt3rRHdPz6JCI/PMen4fyyntROln2xnaOth/tHiULKAS
vK/AHaG3/Sc98m8KLUi6RyPF84ryexyM5oyoY39nZpB7MIu4w7ePK2GiizH8G9j0A+BauRo0SUKv
98+vLfrxO0WObMX9CjM7A1/4N+92IgYKbvqu8cmuVQ297wQDoa+nivTkQgboLndaboR5k2TTt41U
lO/RMMMDFGvxN/RQQbt+vbQoV60fb+ECaEi731gbcUZmghfuQKCQT/WlcpGQhm4IgIgVVug0xM+V
hB+8ICtQrWDl+bN3BcbbPeI1zdUYyMPr7qz59GhZ9hRBniReo7E3AZud3LSGp0G7xDNFjO9ctmGu
W8MsXclTYzC/MKVWmk1zrJH6RWLuOF763CBP0xv9iDIHROnEQyZoS9lDr0GmKHtlxOO8R9AiHmnN
SM5mPdY4lFX2OWDCyRnUgsFDmP7ylM/fncGxRDXVUnKHxegFQPZHuXfYj0JGUI0r4HvNmR7YXcRu
Iwm/rLij7AkiRrozJ9Ls/uS3YfZK4rq71WbJtHZ67Owqxz2siQ04XaChD2D1JGEfTEAYmzcR2bDG
052g35eI74bL3ZOs9OeJWWpekCoHhULJ/PJLGnG41wmsjiOqcMC/DQ1RtgzbhuPefbhsrJ2GUMS9
W4JyYl8eYDQ3sL+RLbVcfq6V5aTiXh+tokIQ4xAEXFgWGWt5l194ojL279gsnn5iGZqMy4qbV024
psXLQFRE1hZvZJrm4tHl/Spz/u10TJFxKNKtgFCtCb1kINWBlfTwkO58nw2loGu+NzMIRiWeulqG
dDCCmAAiBxyCK0VFlnS5iAHOD5t22W3O8AiUPs+duiS/ZroBzQzsoP2Ily1TV7YRH/5tHwceOyj9
YNHXR+ymRHCrnzx5Z8GoElBz/JvrrOphkmZHoo9SaAEa3mDAZmON/KHwmBWmmNe8kN8shLwZSw8I
qSf4a/2NNR7v4WmAR0BKEl9qWIeJtSaZ9/3ORKg/CyTvZwFVgffheYbZ5uUPvxcJ4YHhaLiXhYfb
9G2IB4813gUFc6VZdkH8vdiGx0cB2BSwg5bL+Y77tZiUPfFFhh6aDxqUBmc7Sx9zhAEpcsgXpWXv
/vwPEMhd3l0+Ptve+mlp/oYsIetg60Tn+ZMqJvQQ/p2qvNSD/slS1k5ejoRxli2lAKCZ+TorEazu
PvhUwgfUwVG8iIwgXGSAml6ubq63SY60rI91wndXnDob/lIe4ma48cx8WwCmWa5Vj0i+mnHY8Jc4
QmLUx/Hjdz5DY6/Kt6Mvf0oS1p7es8pD2vZk45xdoZyPH8PGV3HiP8mbd6yol90MRPIW+7Zue+fj
SZdHpXKt2OO+veyJu5wMqnOaHHlWuUuRh/g4ohw5xoIbLPC2kdMsFPpwwS3I8zYaIzhGWH3XUPz4
KzNs0+d/dthi3tjsGi1sZz6yt2Nt0grAkfztUgWu6ccg1Tmkf1PuomTgyv0HBh1bvXIaMc+DKJo6
fGiqiXDWl5pQVvMNLdEi+N7+OuNX984tZwxDXfpIznviAQfp0Po8qu72GzbD7G+asOdhzW4aYeJa
QH6bhYMpayU0igz3O256+hADB7uPZpbgxlSHsQsAasZxNbdPw/aY0eXQo0PgD1KCFzjXlFFmvgqw
qvLzAbgHE/ZE7R6mP3l8VFGi5k+sG0/bv6iDzAYl9eEDJ+NuDJUU5JtFVCTOK1SdAtxxplkvP2HF
Ilds/EQYCOqNm5kqSsW9q14lOdxea0AhTk66vf6mv+IxQmK/qZ/ojmYfcMXApXTJu4NEYCWa3mw5
aJDhiLXnPWhOn2gKmyM39IyUorfNoLki1Ifo8WrNXx9w7YZ421mtBztGtSThXYUTlv6p6Lk/7kr4
WH/WgleTDvoKczc1hBKZwHQqOOm5g0ARCIE6wqBPblQEqe9wCP7hia59n3xIkvLz/B7RzVKihXGn
n/0/Y72Zx04LdW63O/yRDb8ks1gTuX4b8Sy70O2jR8LTLi46CHNfeeh3RPvfoazW0Mr1JyMTulGA
23T+2dNluweXX8cghLaFT3aaXFA7GoSSlqp+Eq9FrCQPDHf7YdeRm/JdujjWdwfNoEG/xADpS/YR
k26c3DkJMwnM8RqwjOW/UBg2fajT5V9pOwGPQurPzaSJ6rccZdvqmjuNrHL58BrKuQ4N91N9gumc
PfOxToyGzaFMfUW2nU3GPOVBPd2mqPUJ07o3IbFGgb50WZlNOSisfsNtGe6XHHN+QLpIeZ5uN/X+
fX4rGDQWZxFetGKfBsBt5EiX5kHCz+XJPysGWyU6+3jxZaZSa62h2NgzV19u4lZ93C2vdQZIpSKQ
xkupUuFP4czCMg8QYW87596ELAOXRZWQChme7eEv1oh3hOnm1Mxw/bhTSycZnwl2Kj0uEdiTkfNH
tBzZNkw2NqMdoWZaeJoDkm1Dxj/h7pcBBRK+meRNH/muW12t8DDWtVP6bCPIyFibBkraePp48TMQ
7oKn4jIqHAkb4RsV+lg/2Hj14Xdptk7aZjK8qc/6CazfEPwWAK05JiMfD5xy+pxMQU2oOLKCge+d
MDcvR48zarJBodlw41pmoEuwsHN7G796j8wN/UNnvaRU0pxfYIEXs1PDsSM9FyM42ukne/86i0NH
xkdNm21mgEUDbG2KsScdxr65mLObZwZUJIM3wx4IBnVdjc9H4DYpTS+/LT+F/arpPg6i5awsuXBS
lxgTXqu5qNsFkG5emMSMC5OodjOG6u4osHhT10HloSimuDu259U35utb/8oyUOaiznjZ0biFrPPm
rTnHxjQGjQ2L7at2s+JuGlFeaAeSkFcuZN3hYM/nzmmBf5qmETSK1Qpnts/zNh6JIccm1CPOhh6C
hsWdepfHq7dw66hbVrnu3Bo7S8r/oxC0Ic11G94WmKgLHIIsqKpJUNXQ+chdzLJowEXDQZaNtCIU
UbxuYrF2K5AzDUuTH87tgQysbcuCBolV18jYoo2HTpovwllQmkKB3n9hFBu/8mFhopAYPrWIx9MI
j7XUCRQicyK9xp4z6MOx9DsYSBrFxf89NQxbYct8JTonr30bH8XGe7EFZQWDEfOeOHnOqEJ63PK0
0gYZZzkxCSLd34ej73fsxdiQdnb76v2HHE2sWaICAgq4b19A9UH6BhGotWI2w24m+nhYu8Nfp2eo
qMWr5I98i2HvTbwMp9MDSAjViYsdQilhTbDsaPZJpdKLaftj1o9Vvv8xNVHnH6hOtfZ3nIXmG/FQ
lNnM+JFaqMNzRX+vIVFngjAiPMfCOT866IcTA3Y8zM16RGaM/EyMkYqXwy/7XVjsf9rnEnuo96aT
c0T+X6bHwMAVdgFp5cJBTgcHV9oMqzFjUnl/2eWIBdYKFTaHwhvv6lfKd1eRdATP9/L1L9BlAKvF
1HbeBZvoA/XsJ+2A+GfZ5jE8uaX17YRti75yqnxyFQj1uk7cg/sOSAe4gHEDFNHzqCI/FHV+K79d
CigIlpqDMlYMiWJWi6yHa/K0arnfGBGKGnkGUE03wvHNc6oxrKT6CPJgMPh+Q4ADRtAKGKlWYkK5
cnA/tXihen4nUI+e4+Pknuxc7TFEmOot8osGAZ3HQimZaN4w9fqQZHIi7melVaeXDxmsHEr1PMZD
rGvs7ooJONtJIE4S083QgYmIuZpJZ1qw/em5/lRiZQFCVJsfr7oGWXg7BSAaEDrEI5TtWvPZCIJE
X+MKsmuTv6qgSLR30fkW34P64EscBpQbOhmAdRrvWInG9B/cshKdz6yc1/emhH0yocVUJXYNonvw
hpruPyBItsbzFm08mO02LqrQSjT6dyOp/s3G3BqcdaZ26VXROQByz4P39UXrFgDShIWhVII8Vts5
RIJDbhTgVVB3YUuSnYxVIG3uQmxpmo0hBVYtYAufPbMKpwylebMxEQgqHkHxf3xKhD7BGF3jZ/3r
96NZ4wT6U2T+tjmZNfQmotTMHDrts+WIpfH9LhaV/51Vn03AkOoh0nRVXyTtvHmGJdiLPAj/9/1E
13FJ6/EMq9ff+r3Q5RKZ6H/HGpb/ucfmo6pe+PmmYWPosrZpzRnPVpi7awhP2Z+khWjJhlfWhXqO
IpIBd3upv8wX9mcI0pUGcKNvKprxIulBOSS/rwGlxsTyoJrq0aBQspzIG3eSZzTr65kP6tsRPcY5
mEbCA5hugHtsyxFhq+25uvL9PyRo3uDKVNZnedX1JvrLxcIXIAg33fF6FkvICr039eaD28gSkIKV
aHlyK2WWIxRf6tPg4v/xPPxnKTdAIq34u8Ch1sbQ9qvQaiyNPuFsZhOpi3xTAEOhqfedzawozvos
bjXFUauKxYDubU7QqN/ITjLlAHPaA3dp0DPeKNgITB8PSuRA3CMo7MBd2/Ti/DNvsfAI5pduSiK6
Q8sG0Hw3CKk0e4sOYpDWis1W4mq7rjErOD+9Of+T20Vj41Q0f8Vwhw8XAbQZBs68iNG0O8NvIdjb
7ZxVPReLqieqJKgpGQ16KMtJxStkliWj+jXaiGWyhUmZMESiRs2/oFnEcv64pSuF9tjyXJKOtENu
VzwOiIKcA9pNXx+Yho1jOkskvVe/N358LbQOvnD7HI7ZJv/JYDP0BFs6rkpL0HahdedO842hSn0x
2EYc8VzyCMnyw7CGVveJ5sPCrXit3fAh/fYPtCA9ld2jwz2xAICLjYM62MR6uHqRy82p2FdhA6PP
MYsSnroEwFBs/N1mQJ4nLyie+QKZZ1p79LldnEamdukllkQD/dm1J6mwQ6xtnQMT1cSFoEQs0j/R
KJmNSM80C/kHCTAfqOkNcSAQ8+RyfFHRKBPflS8E58t+IjZATCJuORh07zYXqDOhfjCRlD41fAQj
pdbVezi/AxaHaXhL+D79aPA5X+Vv43RPlQYA8zRznKguTO1XhA2e21J12llX7xoD0r6FC9FCKeSF
b4tn2neaDQuPkJVGFAky95siv6nkj46Ker031rMRsKDvgaTJpPTcI/ObBqkE2EvElu1pDtFZZkc0
mZ+7ZDIR+HrPhbIVEF/4Qmyo5eruYdJ56qEMGG1ZfnrKlap6G0jWLCTI19mlXWRZuTWjCiDukBie
tSELyzVaM3zXYglp670gzkU9ktS+mR3bixJpBYlHS6AowkxL1viuS9z+KSMBG6L2rgQ9X3BuPavY
E4BOq6wVJboDAhVgKsR1ibqAk8Ior0rPB5oPWABK5V9uo12G9/uMbDTIwJ0aUEanu+Od1Zj1lXMS
gukgYW/YIUBinFFLUw1CQFScNCWRrcB7tRMQ1zCn7JDsI+OIc6rmdg59u5Y7ODsNwk8eC02ZnXlX
jkVLRL7E1AYwqYhQJBvb3DqFf/QcuUMsKQwgwSYjQQNgy9B3rsGZYsF89J0VkKoefy+iZ+oca/5S
5p6fes5yTyxfposrjrCUpuTYdLjfFzQCQdS1dzw293fioBJ6Ht4fA+PWH/MJC19K2lOoRkm9Yf5h
RoceCbZkPA/zlNGpvft4y+dkemm3PTEFTHpMXkwapxAGLzC4olZBWUQRwLer1UQ8FzxXn0UplGAO
7Xpn1DqvTUNBhGZ8eTUT82cmNij63HM0bcv7vTKUGoSj5nVtuI7DEIBNeyWOWkLZuPT7A4hwaUgc
3iFxrlmFbqO8G4WVtQvpmeEUZwjLGiqLdhcxHY3EKZopGxDGB6t9EwgxHr++4Fm3/6/04PWcIL6G
0zIbSiZF8HXaZ6Op5txaNLiYPMVGX1XHRs+jV89irqhLcdOr+zSMBhaWvfNFMYvFosBWFi7u90D3
NSamGTvBJaNd+IRutPKxFNQx0+1i6VBz8dhmbm+fjCgeL+Yur0/tqKIJipIZMqxA0g1k5y8Ixttz
QZ/pqHUyVbh3YrkcBWnJIgRjXAfaxeyAZ3zSCGcUe0SxXVphLLEsLcIFIcKALDx90C7xBi8cUjHW
V0r3bNfv0VjmGrI4Pf6JgsjVqX2chZHJRIUMUhaRt6xaQDqNbQlkYCLp6ucgjKtmS/tI4h8lGaLk
dx0gZ3Pu2hb1OxqPreXgkeWR6vD7AxLyFXVH9i9dYQTLPRVjT8bC5TeD7tbjezylmIOPIAz5yRCU
yewsvvEGTTNMWAG8cj+HdItnadqbPntcPdHEfN9sNI94+WiXBVNrR3xb33LF29gxBG5F0MIej5UR
zYaipzj6sHVEKEuGbs3WLHPP2FKB4vhZj8vsUjpyCZIlfQ00WlqqvZbqsGkIXdib45Ki81Cd1NTP
gKlCaxxya3/vghgc+FilK5HhzAom+34j0YH2HSlmukl/Ba4buGhX+EIZTu9w6fLumR/TSk95m0qs
wTPCbw378tUYnImgxdtWQ5nhWiTXh5YWao6gQDlQsZAbaSfujGxgnSf2f8kOFaFH01TKL7QCjPS7
Yo4y6gfFRL54GV62uXvg+57KSScHLkTT0CejQeyzqY2g50KB1D4KPp+//zlvFimb3IzWpAW8YRRI
CvtTHpqrUknGhT9MPORjE/ldIkx3hQYDzbmMsSTo8CYvIlopfGS3EWpbMq0lYW5AstbqHYbimNIB
md9gimlN0jGol9p0GA4NB2Pa2Uv/MRzjwfyhfo0P3EVq6FDRj2Zs2IH2c/DjlqwJiNOPgV72I/AX
mg+i7inrI7qVbtgVl3jaBDGukSf9+8GdIg11ccgVtJfh9G48fWdCFUTwEftJTbziOpX/ahQAFMUG
sHWd6v+2IZnWB00oDhH27GpRJ34aqMwpZcMOJjMZxA/2zCBzo8xnCGedGsBZ7JtkUvs/sNqzhlRK
pxVKUE7JVqhDcRADa8wp9QfkTHsYs4/OASWtqxTEAznnhk1Jd82OFtQD0W902gBYsh/TNSYINFrr
W7VsCD1weQrJLGce3PxdumFGLKJ5DY6GrqKsJkVSaXTJETQrbdcM0dvJH7+nDQoJq5VwOMsa17s7
k/cHQggjUFDwSY9VMky3bDtfa5gwxG+x/Z8SsmV3ekDx2VXe/2At1UrRq8AaIZXk26antV3MibLS
Suk6/v9SSagAdOgw5kXZiyemQBvN7hj/EHMPzolFoYcICRuIQgpHGNrTvlD2OD0Xbf6qASLwENCY
fVKg6seYK8F27zsqlRU8nVaDPysfjOzNmmffeslTvA2VyWmle0gi1CE3kDvW5Hraxp4F3lYHlkOm
kvAJ0lbkI2d/1ZZwwlOWvH+tWBL77TVX2qSMQAhi+UGlj3290A3xUBSTvAGS/vF9wr9zeTPERbmV
Rrbnde3VbIEHf7DOyRexpLioukGsYNFJV7L8XRbgivOdgIL0OmsSeATe/7MaNxuxfu8NpZfbYQZo
hq0NGEUmPxbXyxAvSUWn4OAKtSe1qCfa+uE4BUWUQWKcjhKMKQaGss+wGpcGfkjKf2ho1fShwsBd
eUkhL/6llAS169KWnOyFipivXH+yZLKRqB01re0eD/IQYSlpjti1wPqRqe/mtVumxU2wNUEt8saH
/+ef/OGWOic9gRiQpPBqUUvS1+r5zIap/22AtaVF+srHOOnrK7XmMWYFkqxM8Dgc1Sv8je8NaKUT
yGjNnVAdhhlumIeEIMaIOl8GAM7UvmhJN/lMgo8EWzz8qtcxPxIJVjxGnGO5Txa7VPX+xDhKsg63
LUr8F9wLGHPHrOlqAU0dujfD4PQ4FidTjDrlb2Z9ql/A3TmDtw7dcGs/CHWvIlFn7jxn6+9KqgVi
ULArd2Ur45qW9CH2UJneyTOT6fqbCPih55rAC+EYixYwDqh1CHmGCTUpVgVffY64TCqg8m+lEhN4
xxEqCirJrIPOh1+oapRpRDEjhZ8rLX7tqIaKET681QvVcUb+hS4R+1i1NqGdWyhiOPtxnMazbEip
TUV03tGWeweshAHTvAtQqJhedzP1syTyFVvChNqfb9jlDdSKm9mSq5gIOJhvY1zo/pUrBhnz6Nxx
4DzEL4UatU3GQifjS+Ze7kYCDNNYpr1WRMBgGC5eXs8HXqOoZ+JT1KghXpeKvd39udLh9ETmKNMM
UsC+4mYBbLAdkgAkCzI37oXv8jWkWUiYwaKP9pfSYSwnq+ftAKoCQOXFK0iyo4rtNNAZ++vqOddA
TAcRcnpVMH/rqtFbV0PR/iDVGvRmf9w263Kdlgsmpk8EZsIT/E3y7/hN5UmEQQpkw6FRJdCAaY1m
WQWtSRC6Z3FRWOWRVOAr+W6NDn1Sl9eiuElcyr5pkQKWs7XpDwzWqfJ1YY7mtpIX1JYDQS4oHshr
DWMqTtTWCe86Ru3+qlCvM5q41hKPB1rFjbdMrLDDiCz91IG6O5luAZOvGLsxAwJ/Y7a6EDTWGL4c
USBaor2NJD54PBVR7ntA3KNPKSZd9CqSlrCqye2x3PN5+oGtma1a1PdR96RBBnTGZjsl1yIJePtg
J52cnJK2+QZZ3KPkyGxvRmaAwH+7tx+SO74nnb3znMVbRLPtAQMcbNhx0l5iDLK/KjSeg/W2Aq3I
mrU5X+WGDBqi3GukJoj+yxleBCAiPtWFCqgKCCTiY4PL8siRORrkkjIr3knJDmrnqlWpxNa4nOxk
v3jkbH6iymolertFSTyVDyAIqQZCL6tBkU02oEAjCZU22BLfj4gazt0uHjqLG1IocN1NozRmekLA
UkO+Fxz+KI1JbGjGoS3NDV5VGE2J700NEyw9fY9Cfo6bkdIO58nCe3SLl+GatDBC9+J8jxXACUw7
FeZrzv0Tlj6OajPrGq35ZoqDa23lMSXbL/RpeELkFDwA3Jnv5ppi2lTsEvpDDVhJ8zgfpitaL2cc
PlVNbB+JEqLEqHnuKUIo30yWJs5QHUwOs4uyRd2WBxibhemSX36NBGF+vTpiXSwSo00ort6cePw5
RKFIrfwcP5jZzH5macfEHkosVi2iOmUftfgPBOCUQO9abEtWcU4G6afn9rcVjpVeb+N0zRf2+BLM
t2D/2JeaKIJ+Jn9nyHBXxxm8WzLHf4hqx+JdNukZll55vq0XhnZE9mE/7n5Gwi2VgBCGWsPohxbt
6XACfNXp8jBq5+FzDcDAPt7TizkGrhcPJY1QPbFoBTwAES454d7P5JsaOfyl7eZkKds7xQ7GqJI1
pNad54JSHd866/2AN5H0761IP2x1pvVc3dEBO7C4fbtkYBwcIIUuJXrIvJpvyQbyWHHMp/Zuo3Uo
DoobnKWlJiCGAaCNK/ZTE9jpliocF2yomkM1yNWOWDIxY5C6rBPuGfrA9AXYCJS1lAemmlgvf5wM
lojpFiSZ+GCPxibCPjQnY1vBKJqyIqzkUYN44gy15W5jlaWjiccODJUgQ7ze3MwBU2Km8D1AYEu6
68bveyEiuTsL7hSk+AO7ulyF3ZJEB4F2LpZc2og4E1gmMhSiTs9VMbce78FNHHKbRU1ilFQeBTxJ
4/yWXmGWBUJB80DJ79vaTVn8/EZyQQDEekqCksNhPlvu6ncK3siAuNGFKgtqPOaE4wJ/nHA/KM6L
xKRAXMdAQHNpVBKtaRBFqygJZeuIKDuOQJXyY3uOvHsezvgG8noR02MG+2ZJlShqOnxcmUVw83Ib
g86ARTe/uKqBlx08/r3NoDIjnI/hlVBvKyoUOtGdCTSECmZQ8MU+dxEZbWAaA/rVorp8IX7d8Vnl
/u4Ciz5h+mO4LWGRmgMAMcjFTXYVTTXcwKa5ahWndFVHCcPwbj5yUWI0IWaIU8mYhY2pF4yC+lN7
WTP2CiIMFYqbvFX6/UbX3o9HdTzUcqEXiCfD1jttWFI845aJ+KCo/JdG2NemuC8iIJxNfRXckY3H
CuuDPxLOH6jpFZEl+79I5xGOSBtPj0UfGFrqSy6BjKf3wyBLIQOcEhgkrEAzjH0D3OqPjwtzrgd5
/Q/vdqDSvvmpGHtodNrAt49X4DL3qzh/Q6mVBw7D0mdzwZXJUp1OmLlGKlTJ6K2W5slzcuhmsz3F
THnez4YnmyXc8k6ySA5K/VpdTgiZ93pmdT7siK4rauCEtDZwACEaJy7F4vJORDtJxVBdi03h0Img
27VAVcp9RbZ4QYzYwowQubTy8r3w0Na6eswrLLK86Xs5bdGHNnbOFqBs7lazF+mFxuzn55eNKMMk
icswgVYHPOh+1pGuHh8/qWXcVCxH7FOZfkRsO//N1/mU6ll/evWdma7RmOhI7hCwNU7djTVYZd/M
m92O3BrE6nXkcIVcqUwEMUT8WR4hqj+SR5M1ylcKOOtBmkFJ5RO0n29uDgPbaQgGdQP5BnfMXxs3
aWVQX9DRZr4+RcqAbS7QvfoKcHxYVDtv2/APMK0J4B79C1a5RFvzCAxpeAhH4Tzd140xw4N4LjcC
9lXI73XP5YoH3V6INif2sdxNPAyBdI/VwBJfxjnlmyo/uUI0Zz7cKqbre8RcOPnB70EOJuLgwQRS
KwuIfYOnuQHZDpMJInDhEY9dr5dS0BOkkGjgthwh7MAfph0NysnFU7Jd1REGSoZCKkZzSL8fhOou
IW/44L3thy2syYSuwWY7CkBaoKzNH4PYKQwQOQw7k7CHZwnCKN579Wp2vIXnMFjc52tVlIdUaDnh
FUK2ai+2uVKo9jqmLcVgkyGKbS8gADfGNNy7Cxg6YfFZ3aaV5Jqp2j50B7JQhVhnYy0LCmxk2xf1
YiVYPyIhaXqsKKU3Kw9hY9oYdExhzUMS6BUUPGc6e9y+mS0DuQI/uXqsL4Wf5uQm1K9fxUwQD4Dc
9clSjVtDXNfYUTlx40I7Jstf9IK7ZJwXkN+wmnL72w2tAp0xEnw4EiTO8OtPe+dmST5zQsW7r0YF
zWoluj+C5oEvAgR2WL316s5H0aksMW0QBLxnlHn6io7YcMgHKQtgdzXTv1k1o7BZc93sm+A0gp4P
UawsIqitrtnML6f9lM6OAZWuo+Lwv8Z8i2nUisZ+/CEQQyg6Or7fxTj0T4aYdxmE0VWR4cWaTmx/
bWtcFtSCKWtYalVhqqiWwbagfNXb7SZtPp4hJmtFbagkdNUSjuKIfwIT8d6I5pz7iE8+vpeDs047
xeULnfntUyi1dyvs48rnnxB5SLmqoGFd8Ihh87KQkec20c2dYWAziNJ6vg3OEzusfe/+UvECV1Lx
Z38Nm13sSNmsKrMIXuxBBHQh8vr6ZXLglqsu+wijn+8CiVR4dYeAklMzs26zKebZ+YmGNfQEaw3S
D399cuFSAeMw2NhrtA3sZoIMYlyhr0dygEHCralfOo+ojc3xz1MGeuh4E8jxk4XRHGehLmH1RRom
b1e2ah5FJ7heHLHQlcr9sC0dTk8RI32hXvVuXOQ/0Ge45UBqIssMoGYeQQYOWBqslOJ3ZaR9hhb+
xF5UVeBQVtRxAZXVk5KpGxPwG8/fpkBURrZdQMoz+7VUAXFxeAF6lvSzf4kiljc1H4SnVt/O/0FO
G7guNR3y/aDSu+BDbtJERABt4pEovSPm9wB+G5mbyO4u2Nc6Y9vs+NtblTCvDrrF8H4laHGVmVXy
+KZTa9lozxPsa/g96utBtxDIprY4ryjGIKCMf8gLQcrtCOuJ0Eiqe1F1d2ktVWRJULWmUoNQ+SEb
7xtgVjgTiQ/4yjUyg66ElYPVRZT+0KopBrDNeWrlRPqEPn09ycjgkBeSNl5IcIDmVvSsQmfE40o4
AYBvvhRppE3QZxiA5pHDQFMc9JMjJzcKgqJtgYBzJevC83rkWtZJG4BmJVuZi8J8Qu9vCw/Tvtb6
0xKxvLhbnvEJDaoheV9AUjl86QDfrZ3BPKbwG/FG2ueiHGicu/pgGBlucAl4eEXzMgN3B7M2JYGz
txcWJ6JvhDkwmUCSFCfk3+WZvbvQ/snQuA1Pjbn71f8K24073VpRb+EFdODyE3YqUBoqpdyrr7Jp
EZGQN5tyMR6wsL6PnaxVb2ekhehbUkU0jL8OXCp8Gpe/uYqYtXiHrruHGfmuwKCExFdQpXcwwDlX
/9yISKLhLWsktJIvxAPxdWoafc0NVqE4z0wraKshSCIcWphZFw1i31fwWO/nwgz2hwSjlFwLl3lb
OyVEfif+hYwlpEHSq9DLe4HIZeHaXOk0XgYTsUueVzSSj+Pws6ICXmF45FnBXXZ4/Dil7pK23V2e
DajNrAZRWLDmDpPsAWlEoJIhI13j3vf1sRn2mZFsStnZyERamJFQIRJOiPrmgNKSP8/5tFqamFxj
CaJXVDPByqaYZ0PtFGgzPx6W6KrzWFfCYS452jmpit7NHZN9WXgjFbE+WUgeJeub8vQOlHHl+rR1
0GaoU+lecKOaSXhVfnCAVx6908n2W40N6kFVwRHk4xSizsQs/KJ3+oF/dWKHgu/QkpE9+DG0PGT1
PXkIODluBz1PJZOdE6XTk/xgeqX6HQswvZ+Bf8VZsJb2tIpfIzgPZYGrBWd2zIdlOYLtAZY3gqgP
D3jNjQFND/DU3Cd6f/puuXb0l0hQPHUSqXSP04FFHmar/R923IwP0Fvb9Px2m/JKYQuZuH13V3/C
pYo0DYKyuXXS0q57uwmepTSklJwNAuYhTJur9f4Oy4kBzjxSqkncyydctjtsXnB2bF3/8rUUYeMG
AbUrM7hNj6/lYg9XZIy8r3Erk9dxOIMG/JG/8u5ADplwuXKBUYDv2PafH3UEsmbevKx+Ntx55821
7qukw0n1jKLZYEMgKqwWTLh/0B8Wu8InCZVcTpN9nJ5dXZZxha4z4RmgP8Sihim4+TNMOEGvngTT
z8Ipp/3Qn8XqzNyiPNm1hS91Ihe680NtZ1Nk4nf3pW2ansT3r3BRxLJ38sPyUdVQdObnRGKWHPsC
QPQJBUhZeUlpHuhtZcbHlTS/mJApSs4/DFWU3C/guBJLjR4I+zyN8ks1dIv1Ns7DCUD4aB7E1Q6H
YSlu4SmuxMUzft9B2yRDJjRV1of/ZCq1zM77aNpf6ajyB/wfikca/VxZMLorJG0dzbXc5vcBEp67
4lHCmtKsqBwti7HN7YTjoCjR+2k/fQvwbb7QaAwzBlnItpQLYM8jq+kBNWFTqqpPqGNMEvdEq1FC
7RqNVZAIBqRjF8xkNlz0rDDNZ4Si2p2eASAW12RtxEzdxyI98wINy2uTT+JINtfn9kEKvZNXUb6e
+zKmZtRYjGRtlGyRri1yYjpK6Cikh4PWcnOqlJR302dd+egWtjykDVKmV5DGRajtLaUS//ncBaf6
sOLClNvTmj38Vbot+YKPdyNhaf1mchRPsCpLruzRi8BQrs49B+85lMwHUgWEugqptq9YXD6aufZi
XImKmGw/ek4ee9q63EilpggHzoLwD3BVqn3kk5rsQKkY+JdgYonSONHiMjDEbIpk9kS+7XimDFbm
qeaSe3TWDjHF5x0ihCcdEIm1BJx79byo8GC2BeT+SviSjmyA+QlPuRSqstxS6BOz/RdxOq6MAT5O
k+jgyVNPgT8O8hmJlsfNSB12XqkpJ6UxxT4LP2565Kj7cqvP+TGj5mwogIYvL6go8+34fsP5USm6
GJ10o1EYaLUiOeyQSX1tFT9GetZF2gGgSCOSGrBe+hBCDi/RVYpQKQsSvv+8EhmCLgW6mjBUc5Lf
iIKV3OJq3hSaU84tjrN1/1VW+1vKvFgch9bgiO7GjJycDO5wciwVk1A/x7knQX97RHnckbRwNpWm
dsKQssOTAkN0hRTcYFRYiAhL5eYvtrWGWUFMHsNShzhl9emT7Vfpm466GY87hvz/g6ADBdYHsHHR
y/+3FEabHsQJl6U6T2OBTP2iXBCMF5tUS4z0cVjZxkv2+oqIDIzRKyzaQRkzi9teC+dzyuM4NObn
t8Yx1HsfpVbb3nWXku5ET9mI9ItpvbGKcPTswCNdPB5NGN9y9WJY6l2MOMBabinsJa/q2KRAAV/X
i84OI4LrKGh0O2p3KYrdqcSPgs7qH+F6CAWWy4sMfRXWWL9W/aMLdZZabsZWYL/k78i3cZqceLk+
ao584mj0BAUt4X54+BLahr/LXLeYkiGiq9U6CaWlpVPI2IpUcZ6eZLsEYM9DQ+KCWD6fvYStvspZ
zcuxTGXz2WYuz/EMY3WwJigTIdumlogi0QCpiTHDyZ59FmKTBBDnGtk/zw9akFwXm17c7W+Xy3h4
DrlKEywpgKDAHiAMNrdTrUh23F8j27iQ/SE5Aysyh93zHT8ZrttPY3haKrzIpLMcbklAnu/U1kUX
9wfDnv1mzVcHs/8xmVOn9Gocrs33Hsl5IW6ctxxRAYWBIjby26VVTJmWrB8YH7BY3D7U0D1qq8fD
8UhhmrY7/E7nNRjDDu+HTV60vtzDlz2A7dhdGNibmyYYUnDRiVxRBw2QmBxgHciIvX942fqRe+mO
v3N09JbX+14iAoE860xw6Nf0KZOrDWBSo+CNLwXe99FExskv3mm52GrNQivsoICLpZEC1/fP6FVS
xEpm+5RmETp1NIWeBOzdvV12Qj6sRUGc11avgfdyHx5yWeXUXsUwiSAhWPwnZ2Rz0Jjd4BZ4q+1R
GilgcHIiKvtg/F9zePQGNWaUI3p1XzK2eviqDqROFE3MJI1NepwtBBTjKaUV/dIHq+XWn70B/uvG
BfLUaYUzflt16t8Bgfz9iWhkZ8uH0uZOK5Ym5fbQrFm7f5QTiNvDYKvwSx9gYxsR3WfokMEGcubj
iBbC1cA2pa5378f05VeP0aU2wpmGq299KcqPyq0MK/k3QAcso6z+aWAKlbn0iemUgEq+2v5qwrXm
hYCnljoN1jkRCYmxpbekK+6NoADFbSQpc+Ffwq/aBPnWjN+epP5vu0ObwiuuVxRLAwyOFRjDyR5R
JGQu3kAa12NThFt+fLOI/PlxQWSEw3fEmlTl5MDa4yr58G9G78hsISmE+8VS0jDtSUvY9cF1xYtT
ZlittRxnUwlHMhiM9ITnjk2zt1ICvt9bG+AJNlxPq9nKOvPGhgFsBAZQYJKc6iBju7+z6n7OMZTF
d2mFFKkaE3bHaaXg6e6gq2Q849gtzzwL+EbbT0NLfGGfN6opH0nSoSKz0ptFZO+/nVNMzoh6lPUi
JI08gTDQX1sFFiuznNvVBokJXJ4Fn9iuWN6RETFlzKLc50N6W2WsMc9v4YHzzJQphn5M8a19HC6C
gxwrmLz4nrpBw5dyNfYm1CCOyDcwNZwPO4hXGFnlYSFLroMzng7wAavYlSevcTvybPPCRa+BKaEQ
LijrFPHIvHKboeiOuIqII8PDuZD3ADskUZAzv+iAI+Y2z3uD8pGvXAduSYfdUm1CUe7AljDumrXr
eXpQd/GsJF0SAyaP0PX4wIFyEH+Jv+q0+4U/QcE2bCFaw7aw8ddVeOjKTDMs56kP7DVoIAGAQo1j
uCZC7dYRJfGn/hWzG/AoTrgzqOWzJfJ34vamObcl+GZEQxxRKyXYfXoEn7HWlmtcALYVDj+c9RG5
7M+8UhSvxc6ScJ72haJmUUghDpsdkzeWvLXNu4bpkOfg066NLSViMscKe3v07aiYPGhCZ0musud8
J+A0/G+p9Ar/B33h7KAd4VCG980s9qlAXu2YpGqfNPuX3xOAlz/NWYSSGzQQE6oDiP4zCgxwPI3H
pU2p4KWjDEguQ8hvMUGqzN3/2vRcM6M9GkHfdGp5IEzIa0e60ubexek6KJuPiaN3xlkIOpcSTd19
ItK4HmSmQFu1tfHMLJpWK/Fnt8G0ZetIk7PEMBi+YFCNDUI2F414+lAdOPvMAcr6An1pqnZPdlps
3+rIrP2j7FqM3aZbzohPws6S/SAgh+fEJzeClbG7DSTSekTfYeV6lNRWxYa/r0skAKz0tRRN6YLz
QW+IlOaXMTttceV+zVZ6P38e7sW54/speZuZo/hWQ254T4I4snfo34SzjiYv0YPtDvTGliLXLRKh
BzfJYPkObXL9Pyc314CUjMykKpMfChYmgCFYTBdM6rvJFrL59V4UfE7dN7QwJZe//HNKtH5UGZ9o
fQl30hxl8TCAaZqJ2W3iKkJuYiuZfVDohAmbTzqF8RHOfzbObCfaMPaVHOONqzDNXKBC56L3ShEI
d/6tVueQa6+RHeZ+zqYPu7/t57nvptxGISIBZ5adWTP34Ka6JcmivWk3REQFzU0T3eHzS6ygvqvB
jIdBXQ8qNeogfCxvC45QV+GDd2X8RYcTbg7QwO0GdSXHZSUxjPu0tE2/MQIJDmj6vmhMkQD0BRpf
4uxmX9qVlQbEZ1qQoNAPgo9sqFKC8+MYY711PoPRpwytnQx2upUhwHvXOU08h8x5qClT98rufA5Z
7iQLIu9J/7ggQ0C0rqpC0griI3MdgCYSoXz8wsnb9OFO5xLRKUc+HMa9+L1MPX4xvWVmepueQ6HS
nyqRVMUrO0BSVDDf8ZbBbMhVER5ef8KPg3+ZmC+N0DQvjTXUGjolgfpnQ+zzJ8YhKbz9SSFeQok0
9OucDcyZu4TrTDw8Gendk7PgYctfiCdTi4+e7NS6RVaAWwWt8yEkiXYKobRHgu/+lQrXG4O2e1fL
rdCl9suTRAozh5ugN6/M1rvqHH73iSNPOzd7MnJlVYu4A3xeLHP+JEwTltvCg1UlVFinnlweNTJz
TlHLSS2mmCVcq8NbPuBdXuCAdIOiAgg6HBHByxX0kjGY/GM+WDV0nAS/wGPxrkA7BYTIGjhB+apU
i784DMkAxQSvaQTsBh80kzqwoSQiL4tVlNN1D7b5MBs9rgOvl8ufiuVBYzcYQuxNZUc/SR1+VKZI
23bgWkJY7t6uWYSwnjTM3AwuNmtDnuLvF5QxKWa+0Nc1VKzYvhm+fKXqdt2GADP3iPwxJ55EDUTt
rZ9yhCoPslwovKDXxgxiDmUxCUKb/X8C8D094jpuLnOoO/RrbD1ljP2GOEQeQvqfQunwPhWigWzF
fbTUJnVBYaqaPaQEJaStgBTV3I8nkKcyNVDY4uncsCeZasVpfBEHUYSHM25sVlOqGnt+QTNPySqX
uPOowir5qBhsK0s7Wa2FLRdpfZD6oM//lOmzJM9FIA+BfmZtKxWd8VkIiXa+yHmgY/F/BBXcb/zI
Xf651hmQbad/lQSZYKFOtcecu4afw0owjoNS97FCnqCthTBrQR3nXIKpSA1TZZX9HTBGlAIY7T6h
mlahRQj6/Imby1YzmJ2J9DAxVfTRiru+qC+yLXX2Odb2FSnMAj6ESPh+ggEmrXf2ZaE7L1fZNS4R
BguetDBeX4MEZz2YDYFY3nGYylrE2GFE29UNSpQ0BgkxnPcmwiDfBAmuBDz2gfOVCG6eMQOh8uEF
Di1uH6KIcIYTULiExXRtMlYNLqnOX88JKwqNwm9f7d9DHufohpHNr96eWp9+XWazk6dcrGD74z2h
aic3iv6xa1hH6l7vDyJioplF5s5zyZR9Kj91FanMvRXg/WjgHiEBaSZOg2QQUtU44uo+xVPxB77b
n0/McIpgJ6Y0IrnW84mJvXu7uzK9XdZZ7zhhTGU1/VKeOOqDKN6pjbH29hQnyhm2CVfm2P2xo40K
HwNW4B4Gv2i+o3UaARWcWGZnSBhwMPR/zdXm+2rJUqlFIj6H4wjVx70GE2cH5wGzk49TExWSle1J
LvPlZmI3o41s8F4qwQK1ISsBlXueox0wlVapBqkBHX/0xtBtwq4gRHTRgnGjho1K1w9NdADa0181
a1ZrUlS3Yu14FOvg9anMgqr3YagIrzRH8rMT/SPp4igZ52ixx08U3hc3MF1mHM2QKMXq8aV/2NG8
pQ+4R7t8FXSqfSMokwQ6LcU+03y+o9PC1p6CzEcbD8s3jMSpA11FeTgZKHDTTZ5+YPZ0hpwk8bP5
s81GlouwzN8m/T7umrYNjNOL/AGqu+4Ij5zdel2jr84wvITWViMNGC8n8iAa0YjqGQDvZZoulDcT
qSKy8ymgN1yUORv9ipityTs2GY/vf2pBpZ92i12LGC4JPq1efEXVt0HZ7qFSYjdKS/bg9b58Dq0w
h2JnsSfsgxqse/vgX5JVBtqPrAkbBzMZlyWI6g494KNcy0X0gs0to3aRu2FbZzpfrED1vcD+nL0+
4VYeA/7Z5TkKh0xCRXDInQIJQopMQE/UKrGUVP0Q6DMESFjwaj9Ggg+cxxQG8lfoAyaCAlUP76Lp
UCzQuTPAhq9DJ0l0LYADEL8dDPP4oim7OlO09BKq0cjJaxC5+LRcDWpktigJbP8/D7ZwOG+Ew9nX
/ZWmvez8l7juS0D4TnBRpM32kTaSEfWCRTd9Nxf1LNaY0Hl2DpjGsOY3MotuWKMNe8PJiEolp9XO
t2oodzHulhNRzbIclswW0gjblbRqdIEk+2JrFCWvFxTdf5dC6JB2ZMuCHIehSbp6dDsWRVuyiNqB
KudOjjAeWj/4CFDtII3oeqe+ACKJ4WuwdCT9ytOdYfdCCc4ZuYB2QOcOBsfdKNzijZEfY4dXyIZf
OQHq6ww5nH1mf2aNA90F05bh3oURBOB86Jn1+h0AaVklY+YoJda30ocXLYz31sHpPDxs4qvg7h5d
jLF74x0tGbHlYH7xv8ERLkA8u2Vl9n4hN2hIkY/W5pbyZxfNV0plXbuQ/QncKGgOMi60eqKKuF50
KGPsasFY6nthJ9MBrVo4NvWiPQS6uAqEkgxJZuF9e3I9LV24eGDG5GdaLSdXC5fER7OxmuSsBq5r
0LG9ddH82WNw1/TekryI6QiJW0LKWnmLxDA3EzIWCkGcLOWzml/1W46l1eqPskbRR2wmiXLMntvi
kOB58uRes1JMGUXlK2ifyt3QRl69w8v95RP98FLm+mBi9u6Szja/7M8VQ779P0PLdpZ6GhoVerqt
W+MxvB+UwN5CygayDUiKiKQImaKcGgqOzX9Ihcp9MXyRZMlYRYUfh9SBo5meLrCE9boxDRcVSTSG
HIiYvM9dmx/P22S/dGENbsHWM2xqF4on437j69U2mDGzcIvOc7X/nHqZ5CVNa+gSykwyBSPsknb2
3inB67lVVGDkZi0ZoguKJRKi5/fvWEMVAZY5ZVKcgbTz4av2Mtg84NrAH8HcEd4sQDZ/xnb8W1NE
Q1Ozn02s1YvLp+DA9U3ABQOBtyukuBGsODrW+blzHJ4S1el0whyXztWLtfLprqCpJxCmjcY4tLdb
IaodnCdnEiXmKSrxBiam7008uIIC7PgYKl+3rzOa8FE7/PSEz8F8NnXpSscjMqaUCbmHmPlV8cH1
Jhy2PwIaBW6DJ5x7/gRERnwkhAo5VrQlNYRzHmFctSXAvXkkNEQdDCnl2yLFSbECxsKC1UShRbFh
1MRXhkAgT56LYWnBO6QIiKE2gAkdSYDl+jRAnK7Rh6VjuQF1Y49NrZkIK54ZIN5bnRsymMs+0GO3
6wa7AbNpZANffCRO3i9RMhCr1FvM12UnudTOl4lseQBHf5oCY/tD7NMWygMxTOxdKmfyzXa1zvgT
XmzKA+ABUICHAhb6bH2gnYZYgqga67YM3/XedopmGpeeI4C//nIUlqX9disoDxuPwrsE+S8xM993
isYYcTwZAQcYeMWgDFjJejfjTNsDlHt131XSS9n7S1L1CYZ7ORh5KbOrYHsthTL5sqJ9yr95evAj
hmkskJN8Lkaupn+KD4lndGEQAypL6Z8M+j27Q62MURpR4vSaidwMVjKVzbXseaweHTMz3kmY9lPo
Xs9f2gVmcM9ocW8a/XZc8O5JczijL5vEryQ4f8m9ad8CyGHIiAaE9Bxx9MEM7Pf41xnTN5iYWlng
e4Viu5sss5re6fTyoumh9ppBgqFLyzZkCUH33thBmkqR1J4eWTOMDcNxLNswvWqEt8nUAiG5Bqc8
34mCGJE9KvP1pj1AlC7mOSzBCZ2VReg1tF4x+2KzFTlWDGuwxrEUWZqYGk8Plpmav3FfROzFwZSJ
Vmt9hTxy7L1J4BZm752oEzuj21YQIeVvuktol7j8VXK249DkOR81YdnYtNb9qlE+Q4knqVsmk+BE
rTfT+s+GuYL9O/6LGq8CZ6r3rKti4fmxRy1aCbs0MMWy/S1oGzcoYlGXl45wkyI9tW8cDvIm3LCp
0pJOkLPwUGuqVIYuLdLBQaHky5rKhC1sKBPBdOKXpClwOFWS+d0yK3RWS4SHgfrDE06RcRYNd1y6
5q3RiJNXBvjNy+8R5UQuglMGbiAE6AO5o7EJy1lP8o43ybeeBZIUVX2S8Vj3HHkaHB7OF0r8+oS4
J6NtACbS7HS9oR5oaHXrtTSJ6CAWcpVEgTMSOdNd1XEtAExeBRfVwo8PTIwNY2r7svLNqRhQ0MX6
p1cNxkgVf779TXw6cpiMVIDSDEoekPMQ+OWwjZ1Yw8VfYdLjzQJyM/enDZSmgh2H+VFpCVkEY6T6
GUJctybB/X5Lh/mu8sVnJybuQjAuogYOy0nVKHnkZa38tKbtdz+kbHfMsyKVUnAvk1in6LP2b1O4
sYmmQXHZeGq2vEa3xJnYkyy2sQofI87jQJP3Dlf9ro6FYeWELdH/MhutkkV9j4Pn+7h6JLKFtwBn
UGBT+sECtfJVe3x5eNb2eOqVnfHnggz8NTPw50Df5G7EGIybVxgyvayor/R8nhKEgYpH0KznTIGA
uH/61Jcb+/MdwQYVl7NHJyzop3FJkUoDRnj9dT6VbLoggJntpFplm7kKqm2umKhOsKs9uET/QriX
rN3pcTZLO7ESt1peIpoSpUseNaaCSDhJO6+AqLBsWicdCMNyxgAjKzqOMl8IhriwP44uTjg/GW8H
DOti7H8sqtkKgwMynAhvKGFdgP508OmTLwYmNxZFe/gr0nElKJhUXRVrgu7LS7s02OE9Sy8fCXk0
a6hvnroWZZiAvc6zhicN/J5CpZ9gdSNcRz/KJDPMAvpnoNLgnIsyF3KVwDziCh/ToWqP17k3qHQa
YjzD0HMwirn4S1vWu39vmRqwXprKEILEwpyUm5bjMFXYbPMzdxe6ClFQh0Msvp/4roi5HzlsIkui
oRRb2NqAT1LA3xjW9RAqrDSPZjdc4DSd+fU9+P67wCpuI/Z+clhJLP4OAo1f//24jfU4DCYcZ3eK
pYegbeJtRbi+Dlnx5RasVp6HZp93/xgMxbF45gs8fHNODX0pwspRMAjDrXtWe8b+1IQxVNXIxz5M
wUEcdT7/QWV9eXxg9yNBjxLuycQFmdH+2WjvsV6Ewdw1tNWkeLP6FdpY+TWidfQNRnUF/vQfTzCd
GxhxxKBBgqNOMEP5qnPo8ce9HtbpdA/SS73deHeAnQSZ1QdWcjO7yo9a1qtPDqkm7v3opFbkuwSk
AYY9bsVcXilpuhRDDm1uKz0Yb9axMHTgJiWSP+wIILYs8K9g2oNBE6lOl+WfCm80QO7ykvf/ObBP
sgbZnbm35YfZIDhXDzYRZfUbDvkSxi2NIWPvJjb2s74O+1B/ENCELaHueZwUx1/F9YkVc86zhGST
f3sakI7+x0rncYLEKYxbFTrhtDuY5XL0x4WarIJ2z54gQIR7UzNPka0RhSB0jLnM32sSxS5qMp7p
J3h2laJ8E+6oG8nJvxE1HV8z2jwLzA6Jk9khOScVGUEU99r5t2/rnjO86lstPGz0eFm8A/Yq/Dj8
C1OJD/JJEGaCpvC7HDOblJ0XxYtGi+8m2igGZfWUnZ5h9VEoGiKMx88P72PzQxkxGqSbIf1Up1+f
9Qw+UTQ8lZuoKZO3rurdkcxmBXWOouOOJ4gHKqQfXHt/OhT0OW+fFFN1caD7CUG0JS21VjHpyw6I
87LcMPmWbMGL71CiNlaLWD/wCoaloy/sJxrpMJv9nDlrndBABfQ815UP9+9oMtIrOmYpwvOIF3T3
NOYoxWhUZZN5N5hynuguuxGLDeOMlpPjtuNSW+eY1qsjl1JF+NWPTn5Ku8+RxufMfsWR5+OTqDp/
+8liRR6EH8v63DHmvyLNpbc88bYi7p2kt9PA7fdWtEm3Z7zYqXhPyxFUL/DRp8fM3rxYVhkLZVlc
EdqomB+3fdQCxCwNHPc4NIas08Yc5Vt/f7XG/q69+XHAespNkUYe45qdzPUFERkGhhIBDzH1yivP
IBeWSKBclyBQCGR5jFscLviG91Tw4ZtBF3fiyXuJqAniWs3I1/SuX4O3DqJJiQV1pSx385rKGo8A
jOLCFVGh+5UEKN/WrGM1MPotzwx4k8+7ltCn9hiyMqJ5ueqzXJv6E5CqVqs7Eg4J+yrZrjWGWQRc
1pp1zDBgpkP6uwZWblyZriHSmAUOgwMEnGcTAzA3AODoky7f2GHRK7F98XctPhUgGIhnjr8mZIed
AaJh+7Nm0rcLxJBtGmYGR5/BCG0zDKoKozW08+SjEhs2e+tb/b+UO5sCd0VYRQl3+yao147KsVGr
B3FHK/dd+ig+Wa1ONJ0w53hfVzbkhapmnUHOw/n0YnvxOI9rqSvsh92kKJrQAb40DFG53hMoDYtU
lBkNqjW2FY8NS1UEjnzsa0z/r9bItupeSudG9V3L8y95jqhpE/vdCznTEnymGRUazFNNEdWFEXvt
zej21D/E1f+sE1PkoxV8e7/yCf1YqD/xgmOXaTHtYNoLGETzBW3MALRo+D1Z5mhPvuv9EsLYCdaR
pQ5frEEsuIwjY0ZR9KfleeTkY1lgr3zcLZVH9vtR8tsXJ+07yzu8eWQhvPkZO0mR3U6N3Ax+Y5b9
+YonNJsVggdCLuBhXNIJdbKauIwHfAOiJUivftb/CSeS2JmVcRYUOxkHkCNojiLn9rivqQp+mLsB
76gUOLIV4hT+LJvENnxxJTyzLnghFShJQGjOR0akiCKLxFEXetejAjouvgvu3pVqT7FMKfl2abwG
1Pw5b6QIAsLZSlT+7foA7lKO6lCZBrm1cHpzeT22+0eLyLtXi+Tp+Z9s9B0YBos+FZNJrhAh+n4R
EVVsVs5SKBSsYhD8FAIPD5piSmVqTxEFrEVuRQ9Czx3Pay5aX4hGo+gt7bGJ5ghY7FgBcA4uAnWA
r18nmko4VT+BNkPurTBi2iTEgQRaATZeGvhYsrI4p2VHLaOd9CFCc4eTsAg2/v5jkdq80ohmUwj1
opRcVtYymIXTwrUTUNPRhz+5eztDYHPsTk+MXKIeEhrWAAgpc60BqgHc4APUMW7AdXyziKL1llHY
l2+jgHgiT/C8vAhw+1ieFuP9P0KnJt7GDXnKkmtis3IZpSgP90Penv9GV5Oqqcy0BHfkGbBaQvk4
FmkW4bngWR6MWDqSQRIgBr77iDqv/1QojVw4WTrj5KcaaYuhfIROYPMuUbI48vy/YTB+DK8qu37v
vgsGu4q/ovBup+xf1MnFBOIjC1tv/aeYLDXsC3iLo9eIzX4GYoUue4hRKHrf7m3IzHdRrS+49JN/
u2IQckPbxpKBqJk2tQYtIAAVA2f7QHGI6k9vDUOO2rzqygo7kS7LHReg23ec/dKX0WmrqUsSMHg4
mKql2hhU8jhJmyPg/9Bc+V6ynWTRRi/75vwOyOILMQ0m9g/RNfpYZhEbhj9HjeLXHQOywaykB7yz
uHbQPreijXUmJUZbvwdoKdVXMtSLfYSTo8N293sjpOjfXyHWVLvA5oUtXNoPlQOa/GS6WE0VZR70
7WF0tpDomowSvYa1U1UC6eL+rQwRijgn+zOdO03N61esvNKJbpcsFpch5BmCt+mwRkw2xnVizVL/
3v1C6h+/DDyeg3bvMMAdxrun/j9V9rhpGt31o7lahnpRroQjX0YuPpLvRcba+ZJ8zYAwONmA2eY7
Ho//T6hifeeWani1vu1AJjAxjFMx1fuYtEmcaoL2LhpAuSdyxCHm4H1VF+IDBHAaeUrrJX2MWMRa
eLlRx8J7ye5oVLf90woufkuJBzHbK02TTbgEpJpJTm2cd4Sp+xEpbRGmNPKcEZIxPhQTdVulj7xW
565hJnuA8Ax14ESXYjFIW85L9qtUzeobkoRtWrLg1Mn7J1+cOUU8sVcHxETrvyjVzDVIGQOGamqL
zgLmJ+JjZCrQLE1iJhAoXPYCQXHfCRqAu3urwVCCmCPBbYUZgD/4EcGu61mMwFHUtl1DAS/elxri
vAEA/kCSVBXF60LlQ38+ZBGfkpAgvrPZrcwyNJD5K1fejco9l2ovI6oUelTvdMkZBnwDwLiPFXpF
8JTd1Wvmu7DClFXXUoSu8WE+INNzbG6/WmyHBdpmb9sMzGBo69fCGZFCiNq4FtTRMd44H6SLCyNi
B5gOp/HfCgiX6bfwhQqU0n8FQqcih87tylnw3ZBtzQpwOV91SvaR/PNr7r6stTLWmV4GV4vV10Xn
K6n+hgda1qwxuJbwomKQPbOp+hjhf7dDXvdr9re7/W0+lgd/wzp2cSvNtJHc++BlTPi1534TlNRr
UM8X1U3LkI2Ae2ghKIRmheliJQvTI4JadzIdh1gom5krFw5CKP4UxzlkBlWfzeknZf3lBV1m7YqV
hoXrAcW4ISGqJUxM8X50AbInvx15KJOdRY5AZ26hpVUJZMuFABoCpkn1HmJuiBc0jUs4DhZ8yfnS
OoMbSSuuUgrd5/jQQjAsZwvf0wXPvSQ2hBfiCKdhyFMsNUh083JAht3/1KsXJPsULL+rgTP47kE5
Lfhl6nepW4PyQlDsKILfwqJBKfmcZ0lp+uHuKsnKOMX0ZLCSfZWXBdtjfkyM63wBIWy+wDL9O0HP
bjwmLc9GUXZYshoCW6wsJJrDvAdRDrpQ61Rnptk19YRFf9bw7jyhbFCS6NTJHG+x43g95dUtlvri
gCCip6xWVvxldoGPGZOmTRYn9PXdmZHM7E6VtF0y4WuTIyfGgSAVyLJssMNu/mUH4wr8jYiWOngO
+M6lh/csSWrjX6COzvosydc5uHojFFS8rtYbXK0mzGgnqHBtvNpNZUtlh4zcgiqFpj81KtcwmN2g
bd8dh5njTgFdl0UTKeRhVyCkX7F3bgASckwcM2Av81TjApHiLUvP5KDC6uiKzGv3kmK6XGQxL80F
MNr3eK07OXd4gomgF9GEm6pRMSa3w/kQ1tWvrPp+e1KBRloLm/s/o50/EMZhuNgF75uxgOD+iWxR
TkiijOcpGQvsEo+IPRRVjqIXi7+kJMNx/TI0wTHeJ/5AvrpeU4dlrD06LWXbIoLd5d6G+HdlzsV1
XZ8th8M89PfLBgh7uz1buNTnZs57Amro8wJQktR5Rq2JlvPVWOpc0C+0l+RL1v7j9O/2FKui7ZDh
fBOApFwXFfjDFByJvi/N/D3ZpEr5+Dw4HnATHLsVH9MnrMf5zLDoMyTfkqa31m/Hxko/nVpCioEH
q4WjJwLl4prCTa4few1ix/N1RMxLY+KJDG9JupaXP3G/2mjxx3qkIWvD7+r2G9kiN4yIekJJjaiq
r1qsjgcyhLJm6m6iDdVuZ47e/tc/RrkwVuPjWst/BNBFq/4HmVwtEYadbLq+PPHXRS3OFOrrAtEV
N9ILOdF3TzgcA33+wekMH35WbzhRyQUF0ejQMxUfDHkVmIAGi1f2DUyKS4G0EpOZSMj6LO8jnWzN
QKULAA+zAiDEK1NLC5f9LtzUGtt6KwrL6DN2WG13qagkHKE6hzpm+dP+RnfzcqI8EkeGYCExkZ/k
FpOZa7ii1RZa2aJ9S/1Fw66OJUpuLR0pT5CUW1+udK7C1FOtKHJiGa/krjk6m+3jrBtKMD6hN5I6
wUDHn4RORIQ9rBMtGCNZCFxS27K45wYSEQVrArIWX4/OpzKDILFuY0S2N62TLD6m6bvtAXZ45cc1
JIPXgpiE9ugNxh8k5Tc4UmZt5R9VDomKDDGkkj9jyTVa87BPxLl5yij4hu/7FHOKvAWDJyMBKwYI
zsjuzk8vgegMYtOeT0+WAv7zh9tXMGyje9lqRj226zsOAkZmU4i1lgnrq1MktNckf35yLrUPqW4k
Sj3FETm9V11xK57Yc5dggLF1eFBDjsMqw/mrX1mqGHJru13AozVxiexn9xrKf2Xb2sWQ548VJ/5U
bbFFCek/7cABNRjh92x9yc69c4BtcYvHZ8ZPUKywuAttN7VNC+qjBlUY4dwLWf3xALyRfUtAlVbU
/a44CsilAXQjMUvIoNQ1L/mWp0fDhHADQHpRWOuEKvX3PcLAIgq4lRAAvc4nIDtHhcf/c0HbsrLZ
7jeNa1M4bl8pGgeXfdN6eF8z88ukeF3Ly/47eC3c/p5MI8zCHmVUrzy4e0Ft2UJszToRLXeJ8W41
IAWuMyOwgP22xAkTldx6lsHmrUxqMX4hCw0LOuQuYJl/TfBwV0ffCWoQf/Y05PJr5ECsNlHpqkCc
pSl488dnQpLWftXGyAqnb6GCGW5pPkjf8QKDD1nKqyaphqUdjodczWuA4DUC2sPyhghUJfx6oeD3
JmeSrHNSwOU6b1e3a9dwzt3u5Ra/FFLlXbi7dxpiFLm7mFncvhDhCbnXUq84cylhCNSNlGSSNg0y
wEKizkHhwTFS94uL9rhXReQMniRZSV5+2066tn6zkePqXHKOikUKylSlOfkWeP7yj8t439PPrvpf
TqhjFPgCTDHKRV+y2sKbrs6agyGSYsr7UHQaAQa9e/ng499JPHVjS/cn3I95E9aDG6migglSrqs6
MbZNNLE9tgM1SZDSuFrE0nkO707L4FHHPY7OGxUM3qH7Nxus19kIALVfpLE1a0cOMIFZz+AahFo7
Lxl1RtSyuSSaOpucNxgO48kYv/s2QtKN4zN0O1PAI/5QD1vUkGL5Ti/lpE4xTpcbdCCHaY6Iddzp
ZOHVXYxyhdfYlsiHZRsdwxQrJw0TUy8fGU+UIukbLPt+EdWmeXNn0SkFTUQBpfCSHfa+/ox6VY/f
ic7KxG/b0ifSyyhhl+zpayG83IEJZvXu4iQVq/Yfhcdow1rf6DbMXWofB9ir4GdMko/cIAy1q76Z
91g2J17hiEASFhq00Yf7n/PC/1HxIhsr9BCtla4uEdA1dKrIuW8c36DHYBgQXcVfFisUMRAL69Nq
6zsXIKa/XCiTJEAfeWZQTpCpzqkeJIm7fjWdGzoSTdUbsdp/iIw/kFcVi/kDRhdryrAACRddGnG+
Wmmx0dnnaShcVQXd1MSQXDbL0y6Y8bttipq07ZLTzLWQo4zbFTU3UwjlAe3fzJksvE+oa9fjuiNP
UBBjPvo7iplhpG/GnInLx1eoAxH2OPTSIqSDiw22lq5eD9P5gBzNt26WfOOVYRhTVppnjR+aEcqB
rZ9U6FV/dxiigtdoHAqGZlxbsW51LPUk993EJ3wGv7GV3TyYSuFOz7yiuLPErz5U/V3G/hwNBI4G
PGECDG26M6ER7MLU7LEkLF3F8jGWgAKI57EdUOV28m6fYD+J8N69FIkcf3jnFoihxFXUrfTHvw5S
HeopC0TDICnMERSIQe+q/jrIn4lnbaQGD0aqjUHazCT9UgDoc6oSIM2l+x+SaYfkdIGwCxiXj2O8
korV2mqIjLXcFsR0AEVYHfWejviMSRJ/wZ8/IrW3/frY1ir2lw+MMIm1beOhQEseUJdsNVBkYPjc
ghcAsFGcyLTWhCg0As3eZNuORz0XLkLuFzwJk5EQcxtjIt9DecJeZX4gV4Ix8M4KXI66Gi7/OM9s
6pp+52kAWBzecY/085Efh9OndFDHBbOcyDQ8ImhoJRpY3WqoZvMtmaLBklDutKBdPK3/GOI7Qu76
AuOy4fFW+RCTTkdbHkjbUuJRp1U1LAhvbYNuOM4JplsfHaHBlFk/z849QZgYGFFMGsBaHreU0c0e
mHXdloAouA6KsbnvGuhLaFSmTku5irH8iQr50lj/wTH83fd1CnMwd80cSAoK8Q5pMTWx/AFj0rYa
Ks8okQG+b7PYhkMAPq6iXXYx38PWB36PtgteCu2LgmFw7ymTfl7c52tR0ivd+M6DQKygKVfxtDX2
TfCOVWvIcZK5Y8yMJUCji6UAj5zWqcieHHEQJXmWUx/eTr/cIafWLgys4POdnUs9aGP6eWRUxBpl
h7uj9hWjVita/PZ9UIw5IN5zCxZthhvlrtlzMPudMCNQBbhCEkDoaIGyXuwJtbfo2znFhLi/A6FC
cBEj4E3RFhrt9K5Y2QyuhxY55yCFPLshMe1PH9QwpmmUAdwVS4WvMLFzZHjH7qkccAtBUxGx6r4y
YtrfE4rbHYehaHEFdPavWrJO9tothg3PShodGB8FMi8AedoapUKTenSizio/JK0NyOvxh8NjVxav
HyrdfEGjxB/VtrBZXKyfQNCGWQMbFGFBzWoRnV/uKIfk/lffegcxqSFifJZKOOvdWfWWXGnfDsBl
GYMPXJPTLGHppDX5IJJ4i9ihVE+cq0iqDqPdvRplkEcItTlLj8iIIdTzImV2i668IsbEJ9nRHThK
GpPK1aPuBBjMQ+Ra/muOLpJ+0HJ1yiEMnEl6xWbcqeH5rQkbOWpqObyHDcHAbkWmNR/4GhvfBavU
L44ZsYmjisbqunr0uEPTqI/ZfSCyZs3J5LDI9TsDZOIVUEIpWcRkm9lUwpU1Y3jZcsjG0yCztN7P
646m71RLD1B5+ri3oIxQRglhjZlWcU2qvaxlyJEAH8iI8tB5X3Qqk4kwe1W8RbL8Fen3dLA8QdLP
IZ00Zthrc6imba4Kr+q0pocCtP82IsCMWyENO1edSwfbXLNfp1e9am+/6zeykxBw2+vkEP2w07eK
qYkMfZs5KJ08rBez8SzusDt+M1c7qY15aL1sndouvD716AAat4CoaERhq41mOAXAF9znOy9oIiiL
KqNph5j2SaMF+FFr4rsD2QPv9HWLXKzNUzY6KpVJBWyyCCBJXnfyg/MbnTmxTpw0mwxOziweJTLn
9AAuKyVbIEoz8Td1oeBln+SOaVzBsstnFFTsD4SR1V65mAeEg6zY3gOf50zSgexx3RyGYKi+oS4M
x88RtOy1PVBNKiw5WUMEYEKUtLDSxHjpvRFxrWm1EPGDANRyqK+hLHNNrVuDU8AygSFpODX+PVIL
JFstbYNU0zWuemGOHdPV9MDCMFN2+Z//94vI36tjcAT/NtywuydFsZ1Q/L0tXbcuisLyqEVX+SEM
cEe4NK4OLxZef6sLhuvI4GF8b2IUBdg8ta70QcwZJQnKZrzAO8BXkzy7PQlyNGEjet4rVermRICM
anOnHighhhOom1TGzUcP/r/UK0vN4EHKTusqFP6JN0lpIXhh9PmQ2vvBE+nSjTvnRmBG7eSjcBzG
WGJaZe2UbbqCjBXZlxCl8Te5U3x0LnPo46pvE5cVB2lEcj8ebCvno0Lp+OtaGBYcdK45LLEAsr6n
Vwx5zrPs5uAheHDUdUtmV2WPgoCHwbUI8beHI4fF2PyZhhr5s9QcbAbQbmLx/lre8+iZIhywJIgV
mCLHrxT4uRo1xlry84KfAAVdNJ+L6IBlAZRlOFXcQmyIRDLHty+BuzEdZh4lVyX/+f1IEUKKr6QT
8SG9J5SZtyDnDonF2m1AnZFkfOltzrprghnW/noFsb29qTxKoaBoXRViaBB3tqEdtDKp0i0JqhkO
nzakuljT1OisbqJ+GnAP9OBR8l9ecR7P6T8UVUZ4y7g0yA5/ulL05RHZIEQI2GtBetDOjwo/gqmO
wFuyS0CBJvoOMamDGW1dHU7OeOUb1ozrewHkUcWon+jXqIF+gquvn7yUJ2Mr5N/LObM/e93NAdvn
e8SORsBYf5GkDzG4zHM+QFvrRcDIjl0k0wDVH8kGqgF02RxOJ0GL2RaNumzWIHCJv0SJTt6zPEcy
OBuo2pWGbx4JzFa7KhQjKkwzrsPlzZlNM4DcJU4Puv+jvuAPMe4kKuDCdqADeRV3FbdmZwboDBSy
cAqPe9woQA1KuyLxXEAb4k3pcu5vsK7+Fxnl9c3glOyWgvnYeI2dOrrUUQErxmQw4JyAk6tUivtd
SzWjzaQuSL8CLcFCXbqeLI/m2vfM0J+OYX2g9ZPg7sQQTblmG7WsJuM9WuPptNdWcgvXB6pdfKuA
lSyUi7a9qgBeR/JCnhwkBY+xzDBozgsnzIp1JM8A2lPVfaWZ9U5F+CRnnwy6Inhau7NGDUxC5HaL
EAFtL9luroIf89yxk6fPbtGrvum3+C+pNso9jZMpXhut5Ohnwj29hq5MUWFbG9QUtG6+q/d4M+/m
ubnxV6l0BQZylRvb1+/aBzZhOnuXj+feITAwsJtctvYPiNMAntPyzd5R0lj5FLNkSbZ4pUELvDWD
/PmYWysFbxYlMzhHDThGtGjlw7ZZILjCw9T/iY+bEs0HZH01LPAeBERm7Sl4zirsG9P3Dw+zPx7s
MOaBM5qRnnbsPv/wwuQFlZSN+0EQJSIPi3hrk4o45I33uLAwICevWgNz1+ZVwW6Q91M5/XnejpFU
L+3oVUn8c9MjbGc0FQLQ8D4y1KrUW/xHc60PeTDb0dVyLzjfxfrqHaFamZooZ4nebaMZaO/Hu9DN
SrDzYTgqeGW0ZAg9TFSQpaafnTB/kGcNHIjoL+ylGCInWU2/rCftm+g3A3s/bywi3QsdizcpRYSX
n7W4/ilYWdXwuzHWrtnR62F0B5iH/boQINvyJg2iJcmCv3SBD+VR95OPzrfGE+i3jPY7v6o8filt
kw9/XsBYKVbKdoAgMMWkje7zW2Nm6LZ/gJ2356PMZSGjXgLl2NFJPrhW/USA5GH7Zf61GIF0bFcb
0Z6NR+qDrC2fy35wvqxSMQ1HnYRZDMM+v3GwdZ2RFtBrVonuxBltLAoHA3spc8z75CykSVEIa5JK
/jETvjDRmAuK8ol61zbI6/M4s+Tthut6xM2/COKF8EinkW9xnSqgf6MXFuQwhvRAAgB3dL18MD4S
yOyjU1U3x3kaHXLcyIjXPBiE5qjYEwm1slVv/8t86UeVQ07iSDr6hGG/qchE947eRivHzp38T9pT
qpdzOKDeyp9EGHqwsigq7dl+wd2elsq/SH7ulUVqZV5FuUiUqCUc5gVXS90ew4rTFsNg9dFybAdq
gTchlHgMJP8aIaWmeO4iIAq4z43a0MYxSz+BTfNbnYS2DD8R4XLI6ioWinXClvBIJnCAJPtCR0bA
2MZ5ZLV43ANEabfOqobMVxnsbBMu7JZVtnVtcRVS/ITLZOzjL03ocFkCOANAxX/B4lIGmxWMTU/P
yPmZ3pYyrm/gHqhieXOFu+S6MG61KD0sP42XNxkK5lxQHerhz0JPtcIkCStf0036tzVtoJCIMLO3
GeRV5eCSYdW5mIwuPo2k+629T+Dfg1RN1MAQzIceIkg65umbO0ghp0jq+/vQ7SK5VV3iDPjIxokB
CV8OIjRfvwXPvF5W9dzObG9Cvq308pAh7hj0jxHu1PKrO3CsoGvSp0oOWqKvl5mJPZUcJe5chD2F
d8QMxT4spkxIqy+onLFZn8Ki8bJ8TsTsQ5jm8EkBaEp8R9Ru1xqK4TCT60qfPnfPLgnlnz8XbwV+
4zW4KhRaVEfZi7XCxCJYCCKuMXcIsIT9bB9G4poX7EqpA2rcDekLL2OkY/SHzuBBQfRXdn57fRrN
tp9St1TpJp6pTMOBF9klzvQ/dbd+bC5EkVyNYtw7FQuW2VY6ic0CJ1PevyvepxzFZg5CXbIgwe+R
HVJ9SMy6OVKosaIKkwN8yHsgH5W4u8JsLgrRntwwgqevgxvnXpo45WWadV/gCpOEIgP5TUY1U4yd
3Gc9Kv3hXRNQDG8SnDiBHulavvcLEcuQZ5EzQalIoqlf+k3EFvohhFby9KJK+EvQiiS180TXj/tL
ZJG5nuOqY0n1lNxqLX+rlxOpbLIKvBmJU1re/WDwpQsCpI/bP9Ki64qDWQT2p0K1j7Vvw53jnoI/
uBs8DVb4oPiVon2IUZEA3lDgaZj1pZnyiBm6cUi1BrKj3GhXdQOayLfKbAHkwDRUrrQZWeVYF1xF
rnMpgWLxkqbDQWgmUwk9MeHipiq2AJ4PqYMMh5tur2QlXzJT8IE2WMJ83yav/QvmOS7q/XnrBQSu
H3+3sGcay9q9sZA5d50A/9pDn3FoMn7Z5Kmd8kwUow0QQz4uPlSJmKVlb7pVvBF3bhbWy5/skqql
mTZu7HFigs+rqJMd6ZblwpJ12LjngNM2JYGnwWoHyKvzPaOXTXvoQ8iJsHfceWmq9MWGpWcfvn58
dk0cvtXGD7N8HxrWm12Kuv/t6eGgRvOlrJC4XUHwMR/R3//TOlnzNlGnlfsVCrCvZo5MDKHbjoM7
y7/w9/XSJy8G16nwJtgUjiFH9SnYYaaBFaswyEOHv0GfQ2y0zMH9uP5iMyN/8jTSduqOoBDD/ACm
OLwwpLDU0NltUUIVtVpu36UKz+Ywb1nFKO+vtLUXT9e4mWSUyYPnHrFuTpbTkP+Yb/SBVRTBEGWv
Z0pYRakJoEolm8FQiEQxSh4O8R6V9YIbpPOsVK/AlizAcUhyq6vmp10NDbWejEelsSKkImEXOI/E
4ZsXB820uR4LRD/u1o5cT0qBN1a4d4HlZ2jFF5PxMMqr78OIhNSdei3lRpY8e3IAdnt7f8qbBYbJ
5wech0AuAAnPNhIyCfUo68KB/R75PZ48PprHV2zpuv7y1c29JwbyRlsBrP7mHvpu9M/70ZIDUijD
xHWsXBIpbeN/kiXuDeBu3ezpbEPOlEsriosWpstOR6Mc1rKIgvFJvbXkd49WL/Uw9wsqjcB6HlSL
opzrLikQt6XGOYph7V/WpKwLGeagJRVsAM4G1eYspBqtIPRX2UR/bOP6Hj/r2Pi5mejL2A5cjBBM
vJvnimT+gIcrW0ajdj81NCYMqUQT6jgO0gd3XJ2OOQZ790XuRwmZ2VaYfatumKPqV0TGbbnoi4RC
sG1NMeDgT3M9aPbz5P3c6WAeull8FJT79HhPm78s737Hjeh4mWbOzgqPbawcyM0VDmhQN7wNIP5f
BE2ZyqdOj57dG9mrPsFcCSORqwxZr2lk51HUEKd6y9YJ3iL+4dwjHlpS84ZZDzXw/DRosGATfrAO
2yg2xhL0ZceW4ZbWKpY3zexPfrLa5mvJ2TxAuSL/z0HW4457Jw26b8LxnTI3vamVAatJarB1o1p5
q3iodFbU3hjVAhSoTOG2Y9726VnDPnk4XdA35SLqM7EhGOsNWZ49E1JwasyBArIfsuMA6gUatRwh
JPd43myoj0BOiWGF7k1+uZ+vu5W1QFGbCwjoesnRDkjfmyUjXQWb2p7FlfLuhuuTlRUY485AENJa
IdIHenLUTRRcrAV38hQ/sD7PwE4WvbjB/iIMZ7T36Gm6ZU718MI55C4QgUAqMzx+IW5IXaEv3bQI
g5+sWBgdfU+jkT744SnJV6hD8t99F2jEv2y7TwbAL1HqOwU44+Q1aGY+3iGbUCA9v3vpaiT2uP5v
ad359oq1Z0Lt4d+uaYVkN1PrC4d19WAf/C6R0N4tvytyNefirYgvVcz2k7rT7nbZsU5w8HsIBpLX
MS/0gPbSfKyHMGd4heUcJjASXvHnMZ90doHst9Mhvxb2zKnMZhSKYLIUXV7RI87v+zG5mwEuZcjt
Z/tVjyGp8WRfBSvdxZWMvOE48qYRB2tYwx7fejIqZ/v2yFjJj2dTTu6r298Jm1HOteXnaC92tXwN
rP4WQfVl26d9QmxPDizPgGQHdLHtTzkg1Vzxj4r/0bu4EaxZkZCYlxyduJbZbcrRCYCMnEHVn4z7
+NiPE4X2MT1X93fDTXi15s7cQ4vxAX8HjPWxmx/VLNrQ5nSqA1sdj3A0xhHwD7JfSRaNKc7z00++
pibKnlRGpLxTnKWsFxSvvhXc9Sez2oqU6wmzZP669adGbasqYHs69zuGRjfBOnWLkuat2eKzT11w
EB2K0h3d4Utvwp0gWMgUrXW26iuqQ8kNVU8N9x90jJHZUS5a0pgG5xT2iNnD8rW1ZtckX+OiF+Qy
r4IZz+7bXT5p/Y+DNl2y+aejn8D0EslBf6BuFoXyh7FtWBOCXyBgJf5pD43YivX8X+gvNwy+exaZ
f/GZX7AxMdTSTGgRtoL6vfYnL0k7cUtoU8oxBdvHTS+CWF6kWLuM5Eg5brzd31W3Lja1TXN4+Gpc
YeZrSTlTUIk/hHxH/ZQRWxIv0H9q2MPrTb1p6RUeca13Iwpodg8Go27YcZMX6/xkyel41j6tnwOT
YjWIt50948yeaKK+88mdU7pj1ijsn/EYO6xPywJb8Xe0jkNU1OqHW1+oZllXgzGVUo+0CtYFDTdt
mXuAUOLzFEvfICDYXlnVHNuQnxaRr5AHHw4g1fkWrR3gXm5SjGWdUOrHRx2D0V2OgWIsQb+uvpSw
5g2gKWWaj4IAmF/mZhHaYMRciXJBtcxJ6VmulUsVCIWt0tq7xnvM3uuXpkmOhSPa/rP2tU29Jw9l
myOpl1/DnPnKeeAvUzmzqzhiPmaSFxj5z3QHmgfCQyugaabJBi9mL9X6appA6IrUl+PUgSVD3deh
INa3DTx8BzWmZdD+lAuPE/waNtrqQl1rQPxefxJZQcCKxJ03KGty69wk+cKb1kfPZD0zMxv95pVx
O2d1QAS24qudO3smdMf1FWufGkGZSz8wCRpoetG8trbpBR2TDXlVaZl3dSkYpfNfG1R/HWbKh1T2
5YIM6+dx7D/V5DHsz2krUeJ53Nb0TKUcXkqlieMwd3wbDVFOC6C05adCBrJkXcu5+AWBRsMfOv0d
jG/JUVTa4przEqzxScEsguyNUXtWRWTttP2ewYrviXBfX/LbEuHBqjJaiWwvDIx73kxuc1cqHis7
+l/40Wx79LtNyBNcy2gYQr5rd2ls6iYqDoeCUIOq/MSlh0cew3kiiXvuF8d6NjyWEaQfS5F4Dq1L
jyUiIespyIQDQdzzjHv4+tBWTu2Ce2ZP0o5So0YcP9Bc55vS9ARUUYHsNhEoCoTqrQsj4k+qaf11
laOkeckW+IXcucEZdHfWZMF0d6l5maHZT27McGLOoKSBjRBTmmtJrJS1RXtkel2RfhfslnnTbXRm
tbnjeqfy72Fwc6EIDKuPUNgNnIPc63NiX3GoAHsRqixWL78IR2N54FiGWjmXSgX/ZbTZtSA4EwPP
a0E07m2SdZhrhLo6o5TlINLXVzH6eGfTwU+K/CH3zqo7ADwvxB46MmHMlUhfXCaWLCmAYsBo26kn
/akfciUKgSKonsHDaZP2ynYbMqtFdiIfzvzv6S0Id4nSuz47Yb0cy8HgC3aqlCdTgaKFycnDZMd/
wkCD4EKVj60qSNy3sCwyUviYYDKweSanUp6Es9pL6Y3h/IXcuUwhhxba6bVqAfkyUkE09dYkc0kq
uN47UWtBo3eA6h5zOpBmTfCoGWevYGmPx2l1SKlpE9HjCro9BDOnv5hiRqB9Lgcb8r8IgPWmufjh
WFu3uQnNWNnkKBfbiXc8EfqmNyChuxrnQ/naHLzk2XsSGSGDm1hhpMsPrH072jSOAVeIV3AHvT0b
/A0CTHeJ2cNh/P555Ld46hEYdISkmOC8eyGt+xc5e3n7Yvbv41IZXLQpj3xcvLzPZsFWc54wYAnm
MDxDi7oYqzDi1UCD68CEUIlyPKt+85OTedj63CQ1gU1oYLzohiV1ykynPMKaTQS0TV4wwlnGUbji
GCj1heuVN7kvFxU+a95cNB89ZZx5K3TeG3L+rVFeqpr9tUQtsnqYlKmp57zZLB4oHxJXHb9gRBeo
C70eD2xvep//s+2UJsrbSgaBDfOFIpUzu8LUL1pMpPNSh8h2VERrZycDDAk6SGi93hjFFnNnQhix
OvqdV5dK9xLwZvbKikdW46XWDEeQfJPKE3MgLPupVG6OuJOqI2L6kMN1DkVgmUMU2B+5H1jRXE+S
r3/aMp+G8QokdRifVNsvSRK9d6KU2EF51LBC0W/va5mBiNO+lZ16goUB57Z5xHHzRly21CqKuqLQ
HxzPgZbcHEm4rxdsr35FN1Xs7A5l/FXdniV95JaHzYl8HzSAmnStKYzl4WADfHJMGYnFB+fqXuMt
DBtr/YIG3a+Z4/nR3A/VMGlqixZFrCrh7NzEEzTIN04gS9NVGE3PRHSRDfYQEVNxhG3lB+RcCweN
GGYXVtzaUdqHsh+QOZfTBAlwC+P+kag60fn3S7tfZfHfiZ+RdWFLz5vS0i4hGdC+vvDyMkHtmz6+
ycWW2MWtbCQ3XpbfNUalkycA6iGpMuQeNTfs+SOAr5zdAcc5KYb/G3cm+w3SpiqPEv9GQLkHnwi7
TuxU77CstRB5d7WlV6GMn46rB76zyFl/nN/qamRuDJlrWsI/pIaUmDSucmhIZNWXmKkCAk6lyq5y
iZxO87KGbwoSUMxSPNI9wbO6gCgusyQl1THby+cQGd1H3Dk8v1DuXHgB+AtLF7CoFhFN+VgpzAXM
PxQD2Lmv5DPk1sE3wSfHa9EyGWQ6zsA2U8O9usJT8bIIdHyo7+MCQoa587RdlpXL/YfYNEwVzdpy
7WhWwoKd8Yq8QQxDO2n6FfMA6ak0oCZxmoqEa0KpvWam0c3HiN4Jl719WGrrCAa7TvfABeMiAsBB
24geHL3q1x7XZQUHRxy3xGWIIj+okjmNRagP3LMoQoul4P8vkXv/rbYgN19BFWupfo3rCpNMPtlW
YMLQ/oxFT6Cfq4a4eCrUzOCByxISaS+TjXawK+2XZ3LQwFnPCmFjCIh15xOqmzzKCLudpLyNJCNv
uwgaKXhFKHAajg51DfKgWKoZpV/xDLI1g5hPk53ldGhKi0NClPFltGO71r8tg14O3/72k2JRBueW
rud2qZ8xEtYiDKPWzy4FIM5j417pvoqBtpK70zQDdGtdSoKKuSCuleeHmJvYEKmnCHYwBahB8Ftm
akICKqBvxq//SYN5oxJr4jPxTffftx05AIYQANr7bW7fj+yIVt6BmyaZTYtPwm/MF/IukQRXxzW2
5ERRVFbjL/FGweiEHJGf6UH2lSFX+4TGA86ZztoQ4wGgXagKdH8Blaqtix8RSjYAfDhP/JcfVi8N
EywIvjvH/EzzVhZFXEtMTdZMQIeGDks5I2kO424P0LytunXpTpKiv5HXS8MJEt61zkg2TYf/6DOE
jQ94/QP0Bixv6t51qC3R+Epou4ZDGIRtxU0vuNO5g5OgU3Bxds0FUzUHeZolr16utr2tUhzzTOcD
OstkqMAf69WfZC/03of+ow5Mz5MscbAIFpgxptrUPzstdLa+jh4P3FPJjjG9WwhM+bDRfNK2c1SC
wRQWjBOV3EzgOpqdCAQfBQP7bS5CbMNqvaYR+mPtzg7kVIBM4Udsykzz3jqhwPgRekzl3encLE6L
jQ/S5zBKNATM3Xr7/dAnLr+5F3bsn7Tga4XPuWcwitCBxUpNbUMOCED+soVhpCM28ZhrsfU7TAOU
lKsqn6Ukjz4ar8NClTBLER5pKgeeorpU1/HXWo8PZY0JLRIa1CA8ZHIWtn0HpRGaiWvAnjsYyavY
BttSjKpMTfmqCP21TquYjoF0EKlr+XlAvhtHZhttfAOClKuqzby8XcXPcoYQdNpc8+DFblgsvUym
WB4Gchd1u5oChR0C/inUxatk39yG+v23zG4OLb0bXFy3E0jFpaZ0VhBVYVgM4mdc1yRXw9FrXaan
G0QGv1gd/XRPWkFc8oor9eXt8dG+dMTYYOR6W3XrE0S/QdCf3Y2DrR/BrDld/pohwsoRWNtb8zOs
NnEEEsi5xxeN4XpPwrCAUkJhhM8UyX4YbJ5j2TclURsaTYBdLyjeetNQno9PR0P/kFg640S7+mIC
EOsG+DrOgYsLjHnv9vjb63UVKHJ7C+7iMJAvqglEHaffqrMMqQ7zjGSpmTA4JowvARdKMOl5sCCv
+IFCpMBqupUmDhQ9gjSv64JSEt95lDbBLtr7jT7rG19HHi3O/gvZG2qbWbMN1YU1vuJbcwPPGGjz
6EVTLgSC4kg6ICRuM8qp0RRVT84N7b8THZ/xQDFTGGRQaofMD2E40eeAuSeoDB8cW4oWGbsB0Owk
rDNNk6tPuMkrJN42ZIuCUNQeP4NSfU3U3+Q3XeYXMgfU7NFRPeFW0NZaWozuSeLBqwzh+H1AZ6ck
htNnw+xMG8r/KSPYbSEut7EowWxOut/IHDIdH9CJ2dg6ENZyCHFlm6EU+e8wVfM8mZGTyrqhJbbW
sXVTp8MlaeqAnC4UPTRiL1lfhnWhgSkghXrMgIeX1YiYriIajggx63gnBowyUTGBUf5YJ3sfFp6x
//d0jspVaUCxvPtRM8XJnDYtt3vhQdEArZY7ZroSqA7YuXPkHXNnP8WEz/eCx55Ww5JihBvmMa3F
KYvJIQuXUkeYw5C4UQypzhz0Dn5n9rEP8NAvMpgFZv7WsWk/gb3s8GjEOuj/9t/lwFLWBqlS4fsb
fyfnq3wLboBgRNGoWUjUFa/jQ5L6R+2VKt85sBQnRMIqecuFPUgx91xiPKIb3dom7Qnqg8gjlw5G
mrWi2+8Z7F0OcwJ+H9KL/zLoDmQErY/sYfYGYbbqbxkQDbsORG5i39VfZo6yZfMzdb8ttV2cfC9p
XGwbnjZj7KqKHrnOmNnxjspHBoTyC1y3nQjXEEqa20gdtchaqbeamnDAZnmwsT3kZCOwhS+mZDni
+tVDv2CyyJapKBRp6ykM6i3fJAl1QKFiHRAPrpqYToaHf4OeMc/aHthkE8WrAvB8gXkseKewOfhQ
/gT2hG8sAIH3NuDpiJTgqNXtm1Dley7jFwr2KyVG9VpA2xDMRbeOVgSp6TbO41+8x7TEcrmhEeny
44lg/ObxLgJ4ZBRWJjHFbx1jK8QjmFYpFt41DwwSAApmlbfYnwQfwQyi0XAj3j4CQ6WzTCLaDppk
fKKQlk192uPmx6ldGAtiKPglnzpS8AKRdERjwNTATwIyTZxkzXZHn5KxTPPqbLSKch0eiwqQiYgv
b82r6JuYrjRHu3HQPx8cYt6d2m+UJeYhgApRrWRP9oG356QN1BrA2YVvgBG0zPM28q8IAwnv6+Nu
vlQ0pDSXgAOm0Jp6JB88X/xGDQ+YYV4F97DxZmJCknDxzuow8IdC8XzmKc0e19c7kW750Nofq9px
ceRfMu1ajGrXqd4cI94hxozuiwd43qDysfDdqzbgRtkMQsNBldKqCEXW/5LlVZDTjfDRakd8PAVX
6tqvh9ej/82/utQTI/q6y1PtzQ+IGic47pe6ohn683Gg6dUJgIZHpazsEWbbK/aQEBvaiTfDZZSW
3zlvxuoYpIilR5WKSifj7KG21Hf1Z+KZv/ko1tM68e/ok3cwewSBIyYOhOvHdNcL7WHVna+eUDGs
GyXDZqjBLJhENZlxgloelcWHIAnZYRh9po6a3D3F+uJbhBy+DXeDrM0dtx/nJZJeQHd/SpEHEWrh
4tunxI8kYHw1hm/STg9wNHNiyvkvttDeoh0MKg1lZKwr3hJcvw8Zwyh1gJTl2oZg/+6L5s1K/+bZ
+6rtotcPSNGYMxoILBpBWdAPOb2Y+e6dDTfkUv92diqRZIDgZdXNOkwpJj3M2Of1AznloH2UBUG/
pSugu7pQv8hNdAXquJ8AoIfG9ARCqHEbhXcUePeZnhFmSkr0ywTLVAM/bCBO7pc8iyekGxbHQbSv
DiUFxXKV2eLDwZ4UJG9wZVgCm+/Q345xIR9TL7tV97Im4NV+dtS5A+RQXmxokB5IuNZp485/E6eA
YC96BSDgbuKmvGh4DQ/jfSad+BJbHXKncvoyRAfAdpV1GC/jtL0fW2FjxKrPpmwx0QV6tbuuw8Ky
QuyxfiLA07yyb7OwCW8eDvzFkhsbKVD/TllAPAmk9h6fJntYeeFzfbvwIBc02btPIMqubsqMOF80
8TawmkHBbOlgOprTpHMD1LrWIo5c9vkoZqieZNQ7g3Myxg/4g6q0ZScl2QL1UUYG0wys1CYhHHT6
9KKBDyXeKkho0oQMOGw4fpzGFmG2NWiVMjmDIeT1e8Py19XrO1gHS67nbWs2mhoKBFvZzz7Z4rXN
XnvRqCmdwzF2S5KDuaw7w4ITELymeQzyQLcND7TbkESHeWFxvDjZwniFConSeA3zXOzan/tJmdR8
Apooh+77TPi5kMItNT7QfBpEer36h1YRJfkT0s7xf0YhXwcBgo5FAFv23z2nFDySNUvvM3r1jVAV
/ACCwIo9EyFv+DtVgVOdQ/KyuXWDWIjPHRgbghAmDnANxrGESg2B9UmMfADIz6b23BdlTyP+Bukb
2ZTTme4jdOHHBqfr/Jhxni8lkQ89N6b/ngIsUlLjbvUQvJQl4HuQ0dkb0E8ZPLxsCdlIS2qXmvTk
Sjp0xoof5Oujb9+UggGvXXjWDUP43tPFARLka3cs2qFSqvFnxx3zobj5tTy57YZfUDnoK3L7Eqy4
Lp0ho2+kbF0rUfiaGakzVmxrKZyzhDnlwlAaL1BuxqFSfdlfEnORTFWLrbIO1uxPJbHqmDqvNnRV
Fh5xNHW96yR2A638M0fjAsT9lNMH4y37/ue49jaurlHFk2PTE989TLfTFsc0XS5nnrENITzBo6bm
5z0I9UvL2f6snvMHEfAYTNdAkxSnxhAOcEPlD5E0SzU7ZDhhysZR71zpTQF/I+2SFYH4nNJrrAp3
paHmEEKZV4USkDgSRKJxoqY9LxL5VAtYhFpOta1dECPCIWS656BHhySV204RC5CSE0mtQYMiI6y4
gLWs6tWwzAgH4cLDNwZbmYAUMCCO78OiOqrYAberBMt9hW1+cdp8caF4656TUUmEW/FovPXqjgjw
lCYDbmTw3mFFTP94vBoxjdhW677MlP2bGHrAgRuhyyYNVV38tDhhT2jRId+7osjuo03N4dQ0kcnN
MhUd7t32ZgzPVv+Vpi0OV5sgqjCHoaG6frFa2IZ11vp4IsFCx6MW8tf37QV2f1M6jW92G7OFLy97
ZCqqO0JWbUrxbbshhG5FjWchvbxdVaz0fI9u0nPiomm7VntS0Sm7RfDnAqiYW8m2DIHHHfXWcK1Z
E9JJOD9scIF7mWZRBFKswZz2URQlWKi1oEoMs4kTWziXcTLk1oMokByJxaT2pxAOeEtBR9P/0qYc
4FVl7cH1ORlNth3i2rNYfWfmQBreX4j6DSHnU7cxvSwsURK+/4ibgUMJhltKO51epkaJS9oXYANd
HS+k6wFnixsZtfaPbf9/CbXMha/icuv1IFZVK2fAI3d5gthwa1BUNvnvolfrChuWVaMb+E52PRtQ
CHZpNSGnIeqv8Qh15KQxweXkkhgCB9AwLVIL2gYL9m5taA9h0wg9DPMmnJKDbJmc1Ixrry4QExV+
3NIu8sHe/Q770N9HQu0bNnyyqBf5V2jSXMAqYrhdnFLvj+pMKRpneadSi3QhHVuYv2+6boC6L6ho
VglbDJHlMBbZ/7CrY0mrQLbUzum3HKOOcQecAIrJvzqaQ9swOsPyj0VezfP135rbxMMxnoGvY+Wc
lntDW3SIfKDxSXPV5yfw+wrhIYo48I5D+xMnElPMpzkZRrAkltepXFzs3cb84QMwGFbEyGJYTwWx
mVcM+6+UviewPctkQCZrvLA89XPkz/VNAv1TM/MpX1MhU96j23f65DkybcVQVu4ZqYy7ijrBkFqa
ZQr7+vAd2E1FokpCKdPqaPVibiH+WO+h+MOfajWY0vXlpAutUQwczR0FQObtIecL0tFbMSqysRe1
m9sPmV10FfD3Zc5TTk3S1e/phMIYBuEGmzDvbhd+L+wc3z4wyVnZWclRdl8QvHeUymMi+BbQvry/
6uYRHfTctvpSpQ/CJfo7OSM82yZ+gKSXVuLHhX9Nq8Bsz1mBRI+TaIvjy62KiC7EkULAPbQkjMdL
2l7mBCR/gaunTgdaprlQA/SJRqn6Odc7Jjp2fUPn6ZoUbGPx0T7nubno1f4pvNXXvQFU9vzpMgb6
D3BEdqhMKAxdssAWCcYP2qJOkwdUQDuFhtQ5Buy5xS1waMbFO+YN8Pq2BKwQvrDAvb/RD5UYEwck
K1ek8pojOrcRHA8+wy/L2ew31knijp3iE0beUyLY7pLjS3ong/cds5CoNK0waEYEaRBMte+K9jkA
RwPlqOxbpLUOiGS1bh9BTYlTFT6HGN/aTpI7eEvdEd2lVZTiNSi/Zr6qIqTht5+CwMBrKy3zEh0F
WNmXOfEgZdrVwCD9YNPeQgPTkHNyIGTo+/ABaKfAzFA7iXxR6ql9vzTHitZnO0QQy7hlXlsVE9ww
3N/UA+pdfZXLHdzSXb/dKgYtGpeFLT21/KSgEST6/IVOyLp8QcjZQu2zcR2Sf8GNwKw2DuS/SPTq
W5BVBoGEXcBYEygFe4Wv3d/doNvt8yJjzvY1rKLG3jOFfrqp+Hl88TqQUndndlsUq5OT3IP8kkMo
wpK1IIDWf1+AadcPAWLoEOlL9p1CEmBrmKuyZHD0wrO64HEfQP1Pu2dlBgWL6DE/GQMV/+nFH8Ta
qxyHEm+c4xhshCI8hgRpEYKVu2PdR5CIl7zWWjpRGGvBlDkztFN7N5S7V5UpgLDtEd51r9R60XoB
EKdjmFUF0rfiFCVj9CbizQOXmgALit+09o5jDTvo2aCAzZn5KLeAIteUYhmLizezm8T2VbHukagJ
RFUHqBEEqqKTVqIBetoBszDMJDKvfehGHPvLoAhXyKLISSss4WiJVkTFn70PHQMgCJnAaoVV0wbH
xyKvrtBc+2xenH+nBCI5ksLO9fgOWf6i1fELvpZ9IVCI4r35WCGeN6nyABTjvdke9dnqrIef6yCC
uFpFORGkwuYv+NgeO7KGmuxwamnTAmDtsRBzp60ebK/yHX9zgGN9hzYvWQK5u6n9DPqMWnqyx6Sm
XlaqsMMI4zdB+aTnd6nqfSkuYU0QZLrifOtKjegsxbkalN2u8jDZNjPBuUS0/ybXCQLHJ85jeL3R
qyhaYqnBrfAUe0loxvgeGJ4JA7SJj5Q07268JdwZNUgdZ+bYKqMl8GGOiaoeATTojy6xT+9G08kv
PcD4KQyofuO48XURzi2azz5bsBaz/VoZ29hhB2x6TUQoODRpqTOFRrKoRAIwMmVNX0ZtdLEvTpiY
p9Y7sW9kyjkBtUV+1QGWAXPBREpyX7DAYjicuZvxo+1cVMAJkJPAiRdyQEfnGABZcncee79DWRy5
WCGmRVR7FugQNpVu8LP49tToPYq7SZGjLWKIrhsx3nGWMeMl1zgCtFtmEkWPI8qiMKRCdVyuruUw
FJoJz2cGMf/vhUwtVB4khdKXZd6kPrpoB6m3ksOAfjncIGLd/+Vso6naGY3xL0JlgfFwCdc3gXuA
txCSIWDQslJWnFuPKI4LfwsyNp6BP7TXLy5buHs543vg6pfm39QWIb3P+oVmsRYxHn4r0r7puVsB
y/XI64RA5QI8Bhyx3huaZr8a06o4YdaJLGYl6556utWXKp3Fkk/cVCnWlYY9VXmbcdZ3CmrhRXaa
ju2L/68VAb0v7lgqI71sS1nHy8J4gEZ5pWVWcU2NXpA+8JHOE+HRdKnMjoNx6frKF8Jf4iNMaRMZ
/bBpQwwQQ7USFNHd1vD2lndwmw/YIqVW4xaQb2ATJrBUX3twUnRQcNYnQ60I9ivE9+d203G+7u6j
zkEHfhIWOLmXKQ667hy8L0LHlXEvrkx/Dg2wwPECQ3wyhX9ZKb8GCO5mFKZxeYPFu+PdvbH0kl1b
3o0XTGJb3XRA8QNkXTijapQJHwUSbk7ZSH2mcgR0/uGB0KeJoEXsL8lzckpkzWfN2rIwJrDprxgy
FWb8MrRTc+vJ0OWVRmRdXnTGYGcECqlK8UyUEpxB/5lmkZwx28qmKkX2W6z50NAdmOMKvb1mMODy
XqAQ0afXoOJ0qnlEyoIxztIcHhC2Uv1A0CsjiZr5wK2WKDCnAWtuBTxhX2/8tVComtvyaDpjjdEN
uzAvohYWs5CqqvOEVSekeP3Tangzo3HYQ1iQQI9JDRhv8l1yZZ2dmBiDIdOYOQEVAhH1dPPiMdf1
58R2rQfcfvLfsyLD/IemRFtluzwKHylrQmRXFcJVNqUbSug9nj9XNClNrmaOq/Clx/+ARg8CeHcl
difMTKBsAWZKBlDS67QVvIiyaDikZYxauLm7ZH2oVxQyxiBbBwOeSOeRZQ8KTmV8OntCvyYyedMA
1C+3NAQnRBaTIglS8VdsJ8NTZpLZZxaC3ayrvRi/lI9gAmGofbxw8/Wnd589RjxLLm3wmFWA3H0v
/kQhimF+KbT28cTX8bzYAX+53vjJwzRvvRFhCCbwuWDjIuWjkuYTnFXmZ3m53PzXPHIMXZoSZWNs
UeyIYEquad7ptj+p6Z6ItPti9/Ml4rSeoQ3KJ/NmumVJ2DkXX8FAqxD5TSfVfYK2hZiTeQsWm+Ca
lzWcRvhZ/wVjpuMtJMaLPuVBXb48T4LNrA5AUUAyIOKOQfiOz8vNLCJWjEHPD3z3oc2BfgcBjIG1
ACPpcSfq9WPrzwzmJQOhH1FxRMdxzEkEFCGWHs6K62U6+IrLtvYKrSLoejhjFQ32BCVPvXmcRA/h
YJqM6ChERe8/Xp4AVW/rDU5aW2kMlXtPj+iNxctGfmjnKkbzxOADBlX4defy96GRDJnspLRauWKP
shy0LMFn+ROqSZQvM1RU19MbpvKfSG747KW4Ixg+Ij5JSYWeDN3ot+TXbeFS2AchZRZV5gZnmgxG
u2gVNgTCfIcWwLxatFZLbxo7F2KVaSJOU4lTUFpAYUbj4QQFp4jVF4yZRYi3sqWyLyhv2vnTAOmW
xbz85eno3csadDrrwRPMhUG1rl6M/d3LOG/WcbeLPtv4ncxLznx1RNJFgLJs/pOAvq29zx9X5MUf
GGiVp5Oda5k2ouT+bcS2eSB2uBjEA7dSY8SE4RF4DM26ktpNftiTwemeeUZF9CTiy3CQLCP/RCbS
HzwrF4jzd3KrPJWYqNYI2aOWTdz00uZdj32BSfJTR4yEkMTm5kkHf57RW3pb5i4RiUaDfXb+HiDQ
ScEX3Q+QDh85Ui87ur2ra9lKi0W/LApi78iCuGwtChWGmwSoJ0tzqcvITHvy/Hji4jBKQFbtVXOz
DQDmSqSLorPy9nwVNUKuEQ0aJdUfJIJVTX49wMLCjH0vQIOT/22oqed466TvdhMkCqkyL3Ol8hfd
7p93p6j8nUxJgth6xmyRx1kvF4I1mZQh5cS3lIvKxu9MCQRVzvcXvp2nIqdLaSjmwt5+iGB0l19b
6YROD+EBLylTFYupfEA98avzW+3D+efBc/SSomkKyy3b+QeYIeKjNJRQcWJnh1ExqHwxZxRj0Rix
JuSHJ3R/wWpYEhLIKZhWIvtzYkNKrx1yGT/iJ7rErZUBZOPbHS3MaGVDGeudsWW/aJF/nAVhXXrA
34qD/SuaaMA6fB9zV7h8uwncZ03BeHwP/+66Nlslr3ocEGYY5ggLrZqmj500g1VUDvyB8r++WKzg
Pjtudsacg8A5wF7aS4W4E054QuiwWODj18fMOMe4xRg5/Jd6j1TWXDPiOhGP4MfSw6/5o9cjVKhl
iYNhJOmAfWU0q046ncx8CkvOIv6zSvbPb31u4j4Vrrf0BUoFeq9uhF++sZVwBcdOi2L8ffDw5Rfi
uvrD/LV/9DgcaxVur6Hr1HXtegSQrEX2Ri4uNph01bXPTPFV7Z2KJJKnMrFC8MoRslHCxws3/BUX
zbovo3vol/xySWebcbQyzlQzs9IldezY1dBH0q+BJjW671T9uFA+079kAivDzXlurkVnqZGT4O3X
s2r/oi9DlT9c6TDOW5LLGjDAae0y4sFG/qRjjTMR2BbVP2nWZqa4BGAnJPRovmOWOTtjw1bfWunN
kWZA02FxmALvyasFGp2RH3CKAljWC9WVs9KA0Ny3PBqbH4j1+ZuWhYJMdq/ccxAvJAk+Ebj3XKF6
5UTvF3qJ0Iq4y1r4nrsa5VLN8sCxV/XAhT2yGF02VXoHoB/TIPVutCBchA6iko/n/tjttmwqQvdK
I5AqknXgu0JY7OJtzwqXahpR8t5G99dKmvA3AGmDZmoCyhAtEbqupQNuU7Jeyzj+pvaHwuGGCKlq
amGNlPl+ZVA28wx2B9l8Ci+4yTW+Ta4mpkRI6waVZ463HhQkOFO71A+uZIhAl/3QQRviCtkNeT4q
LIYbEAt3IsQ2QijLqFfPEOfqZhnlJLvsedlUKe6Pk1Dp5sUt8HJdOv0F/7ODuTbV1p0SCS0gGnLV
0UnAJcYSJe2lWlwBerXMyA4bJTrqEbYc1TaqUiQXcma6w1d1tuQGgJvXgX57vmAjZvGNQ1GRJDvr
9ecLeF3mOCyTWDKZn7V/oMiJYM+GbDrYaQ/4ONH7eFyOkRmgWlpLDXfyoCgLMSBMR2y162Am5a6/
GrKsFb5eeRgBBIra7AOXA2byLzP+E+NObiRVUCiDicK5/msCJu8PApHjkJ0sd9OvxJg6P7BYG9QE
CCR4fDD8Yo/TbQFJwcH3THBUBDbRId1Nit6PVJMxILHg00y+IJZnPwO/mt9vQ8V3XInBy4CUV4Vk
BeLsEWCASJfjcrhqdmw6+TH2BrIZidqdvJ1KkLKm7B0tLLHij+5GLzvxamKmtOdSs39oUQxwRPYP
6grUnGosPw2mQXnRKvTnPKwzmKsLVOccv+eNhZBmObOtl2uCtCv5vRf+gp1DJOxSJd/7baDJyPVa
b80Z7MZUDOKLOnx2lRzoC+1SpY/HHva1bmL9W1VStQm5Km3UctHFlO+2uocSydeOXqZA8rmFFDlv
KorlvKNxXrLrRTsjGnH/2VRB9Sy6iXEpYKGhThB5jucaT0Om/XyZLj6ql90+Pt1IgKDi66mZXKsF
WG5P2ncw81XN4l9R/7UHPWAw4Jodj/0D2/rMKR9WV6WcS6jUVGjAUvRCq+y3y6ewle2WSA3D00/d
VBwhWriCpIZyMQ8pKr3I9xysf4iv0+5T2P3Xn0tIjAyUOQ8U/vaw0lcZrcGIhFLLh2KDxQbef/Lm
OKGjLWIjsrHHt45cz2m2fx1gW5Ow/xRcPuZxTjN2Ia+1HzlUadIa01j50p6Zjlj0RNWKgHc5hZLE
XvKSse1VA1ghIihYpi/pigOi7cyGpNhjh+Gkfp433Vh10ekhKijniMjYnSsv2sScVjoFARMa5N3L
Asut8HatsV9mSuFkeCQLJmiY7+MceUCVZDUfjb/eZG2g/Z66hWxsik6s/OSoh/luYVY5eAVX5X25
FfEeelGWs/EGuirHyevlwV/wzAAyy/f+0sHjENM4kNpRVm+fu5njTvc3i8OZ7q39zw0mzmULx94X
FOLsLYWArYDoIg+oesvKCoUXLQnFFbHbKojOXS/jlDmHGC206xOUlbMDoeDGah953Wf9aocp2CSV
9ukDkCaNdkfm/4l+XDLMQZFOuhCPkdX+H1/nOXDLMK+I00WODorkkEkCbZFdbUH7hZ8ni84+UFJC
0NogBEQNHQIr/PuRYPReoQKowNY5kEBIe9EQfMo2PTHG2cYeTqXS6LkOPgJFxcrGuRZKCZ/p+172
ICQ1OZvKlr4ErswUxh9BzaL+V6fTjCIWYYp1S+k+xvHyX8da28VKQkMZqwzNpyeFgTlbCeTLe0tt
fDhAe/D+ZBPuFZzC8Rw7RqOz/uva9e49Oyvpe2ss86Cu7ZUCQiWVLuoUNxOL2NAUlRsZqb0FyM7i
6CByo690+i+n54LmFzIOck/iI28s5baCFyynRNaqtniWkOk3pYe8LOtxsGFLRXd6CwOX/qnEYUns
+0xPj8Z9GBX4Vb1v0xXJLFC5uSccRlv7UJU8/4ApLvZLcuukCptRvU4bwCS5BMH9q+n+pqw3TBVT
Ccqa+ByuysoPimageq4MVChOGGeuJiEp+zgW4tGeTIGmz/Xh+Eidk+D+QhN/opGsdKOzD5Vl+eCw
HHKHyKBeeL+jUuJHs5XRu0gyrXnObJ6ViZjyTPktoMgid880d/3AvC2pL6jOiU2YmxnhV6c7WQYv
leiqhreaXKGR4pEvVxg8umsdnFQMNtmiT8qarFCdhRBoMSWhDcXaCZyNOBKvMgEOKF1/lm2nnptf
3gbyUOamYXADH8z6IOV1Hx7LxObP/w1UIbGOsKZPgMACtewZ3ZuR7hx6uKMqkDDHl0XLPQa5QZwB
oK5tOAfsCGzZaxYIzw8h8gG6GRtCALdPcrdPzLsoWfXsAvmTuJQGqtG5pXseNTTrxU8fTSOkuuJ7
sTP88uHk2hnA6FELSEdLZ453MKNS5hDs/mmWqrpL6siRN/paFgamEQFwTZJs0gBIstZwRbpCMGa0
Gh8C8PZcReqdtFxMO0fo7xEr5FJJd9xmvmj/mWcce8TVnJyMM8VtFOiAKvBHerj+BBe+5UbzL/l9
SfxsvhWPJL7SNmCKIH2hTTNFukX2wnBAIu28tXOMsmWYDwBP2Y+Zy2frcnJqYMwi8kl972pOMX3j
l+xp/62eMB4KfvdwwxsAvzYOz9z2/VOxMAsHHio8uKVU9Av5Y8eMLS/qm3cUatvLfEZzBIZTEGx9
lLGmvWb9xx3FwhiK0TlyjF0e/1L4MhJLNWnbF7DKc1CFcyYV6ORPeoBFXhBVU/NqSPHQiy64G7Fz
Y1YM8KY16nFycViCHVEPb+3NrKvK4SY4RHR8naX568DzzDHOmxVoYkCGyhOUUYpQJfvvHxSU7UKS
D+auBXcYsw/Korzd6r6Z3I/1NiwCrW107e/pP7GEeD4wjV61y5nRwAGonNdNxl8qf4J0IPHSOxl2
SgMIWuVpzAm/9YobDmx7e3rY/UauoQcyGr5WxHIpXUGnnSU+0GlAL+lhoxYie9F2IO0wDA6yTrec
2q0SajXqgCAGVt6ZKnVPSULBDU9x6dR96e6VPObTASaMYponsLw82kW0EoRxtb+ioRyggEuN0Fgm
QpNBlcHx+OPuHGQruyKdIPSlcXA/AXamK2np2ok4BVyozzTI3Q5iBVkCTtEi3e8jjgvrUYvuAn0y
1HYUcgqMluv7PkXGZRn32W1xTBJuJu8Y3P0ji5xWP1x/Jo4tPH8wpXGtHJVXWeUlv4dEdsokd73G
j3VhodIVduqsNdkWqb56qrtYJRKPuDvWcvLeaVlEKnALBUt03yEjQAVTmH8OAt3rJdMafAm5vrEB
qAGFPCUiLa0rRi9YZSfBptmt93S3FsbYPOEyVaE3t5eyGw03eiOu27EjMXc3tMCPp6kZwSBkvsWL
tYuBs4wv8SJNDvrXKv8PhmogYPZA3F11fbjA9CtcEB/KWFbsXjlM6IFUPpTz3Tz3x9IKlrdVblEd
SD9iujoJS0R+KwRlW6mXBJAUL9dGv3Q1NwPu6ci4yt/PeBtMKPgt+ueVYD30tWcBjp4b5W8SIsDj
dnhvOt5lWvfDdgtyKmFw+xzc0ccsDMGeDdG1j2zdLw90iK4Ye93AOHGxrpaaUv4aaAX36+yCMgbD
z+W+HNXkaNNSn7GYXzrFajEgmku+F4aNl2g0rph/0zNyv8oKjmc8+WT4LKFKMPD4YWQv+CbfREFD
JFZds85FxaJ4js9meQYwwOUVWQt3z+nvTyf7WxBHxzrqYwkdJtTc18nW5H0dBRDWG+iHewpGmVyq
B89/aH47GYk3JOIVyfarLEB+IzPHGpPipac4GEaiTScSSuabG0Ij7jwleOaGizxRy6WUNe7YnmGf
hPiEb6MO7sKabMr33UFcKnPcBVXMD7Iqd2QDDE7qDYNFSBKMCPLTa4FzrFpYqM39/R4zMKsSLhW8
gV8yLKjvXOoo2L0T1TRUWz+CVM7xpMmcZSthxulquy6qyn/cAbnOkw3SQZT/fw6syD/+PCfYRJ4M
VcOi7TLPo7LECuFA1Su60HlWxLKCHcSj6xe+Cf4m9YfJC7T+imWi/6VPR6Z1BVW43Bgl4vtkykni
pK4jGmkEh0N8slVTfZKHiwjhZyAKp3uk0DNBSsBxI0CwIqE9LBBrjqSMFpmQnD24dRvuOKq6hIoQ
hS6XOfU+AiR4kfjHoCtcuTICbz5n+F1pleXzICQVg1rcYkxnz8RME4jbdcbOTE9QWiQ5sRBtElRX
XCM9FRB/Ll8O2E+i2g/iuzU8o5tEeZ88yROa5fBLHxQ42SG5evE6vYby7H3Y/tMkFT6cCxeT8LDZ
Dji58uYfsqbjgRm9lrEOZvjHLc/tZ3CaojmRavvgQPS2MPtEQ9d+/bphFh0Bogpi77dyOUpauPtx
ro+Wt+owilYGV7qIPgiWrQqhDkOPS0tYgzyJvN5Hq6U7Z5UNsA0qIIvnKYEkjYO4cl9FbIjtrgG3
BeVdYK4OcpO3YD9RTVydts9jUoUzGRBfG5eOjQ20FALN3eBkoNzRtugn3ZPNKk0y+AkfqVi6uJ4C
oeox3MHXnE7Gn0T23OFySxXaYaJXfEI2QtdtldYR2qCBWlHvs9VJ/TZ1Qka5bdVut9/Xck7hOwxf
g6t7jyembuOKJ2Gyea4KD3rfHy/GRlFZJUfocfUdMu/bxCKCFfm3hAqX+okkcRwRNpeS300bGAnx
02hpP0af3wlHTR+QIO4cbzWDsBoK7IQVRlLr3Z15Irjc12CZli1V7t6NdakdfsPMrOn2Fk8gsp5n
M8OltS8U+bLmzBTpZ7QNgY27irOvHzOTBkuDE+TN6uld2Rd+mKbSecK4FHhO3/vI1KqpKJhzyAPQ
X2DRaEbT50014teEq4Lp91K+3j9rP4rQSvmpSycfICZPdXf4nj/WEKsoevHtsOV8oazUAEbhb5HZ
0y/yZ/zON0wEYNO/yql6N/M447HBFMH4qM+KPmRzNReFRenuXpL2G6g+fM12tWQvHEPaCx4Y/ORD
/naRTzv3JC5B2l9qyUjthqVWO+WvdscDlSDrtBQPXglwxEgEEEYJOAyeMsdBdApisVC6YZMCb1xx
5r8rrX24C5CjDl3kMQyE1Jse3rR6UBwQc9FjWUa5XPJwCCAQF5MkvRwOiJajHHip6PwVSeyrl/K3
cJ6m6ukO6IXkerBFc49yrciWU1TPbuGakWt2Ps6k6/++S3zUJQOoYsjiENxG2phcKHb8RdvQdpB2
oFJhK1zZjkcemXchT7A61LKN/Vgx6tw0PH0cFL6fYkm+dDH61Kc+5KAK3R/YcE6xrqILIzY+zb4S
0msopj4gy4Z2ULeDlC04PhmJpq0PRU8FoYonMng3GnsYMpuGvcxY/IxyIsVaYy9aYrSH51Yq8kPo
MD5pmi7EF8QAEpNURvWerc7XGKerhbyWKwHrg4DLaIkSyvdfVkUVOH72zHycpyVHLptCfWzr+HEN
1fna+PxmkynIUDGS+rvhX1FNZl37mzBfmUR+KOeL6R3rHjIEqu9ksqECZDK3sy4IZOLLj/E2Pzh/
RHMjr59ebJhC1wQfVNpE1pJwa6RYVRdVFZMx23GJT9DfZwjkWqRLCwo1XbcKzQCRGCYhrID5GQgO
j9Lvx8byTuDQsX7p3vGrJ6onDOD+ZgoHNM760Nwh4lQBpcE7HJfXbY8LizO0E2ht2K3snA6yiyqB
PEj1P8oANRwvE1ZBZyJveEpC8nC8kOwEVNDmHa7aMghpoJIKsAknR9C5/jMIcbTornvMIqDAE3vu
6IKpkw+IKmw+KXIYddQ+VYpwgueuCAlGcBQO/S5sjuwtX/VMMKhOAYUzJ3unSzJda3futTwiChcp
Sgq5vsyYyIFY8FjPV5OI8w4mRC0EEJL5t3mPTDxSVfUZqloT4aHyYGnDNuM+uT5NI4zgqtDdT4pA
z5PawMEY8cRJt/WrpXLTvg//kFfMKRVUBUl7BaCaVU1mS5gleoD/0Coy4iL8U62liN+eCMgx88ys
InpSaado1EQ4fgeG7FfraOE4R4qTUXf+yX7Q3RcCP2Jruvws7pN2gCJLIh73LlToFHjrBHCgIGCT
jlAiY8op+crZN6H7adaErjgWwGNTqcdstcRkfwuMJk7HAD5AO1PCsjKMdMSJ9EdJttJMZ2VOp5R1
qZhYVlWK/wUtAGVA4gqtAkLjq/B4jagZjaUJ3nGQDSu6XXtXbhZNc0pSDp60qSOs2JXYpzciHK7v
M6GRzxoodPZQlmEHV+3qQ5IZfISYYY7msRvJj/vybuJbjDAvoJXyBpni6lLb0/QCzhE02iCIQXeh
3C/GXUc0mgwkRm9Vpbmc2fN33BGh5sWvP9dWoQqXe8hzKWScXesiTCurJ6G0DGA3e/HXlkatZDiT
0ZTkZnJcpNHBXZEtMkdmFS8D0kUGCcrrhlRqF+UHtl8Up73j4/uyKr1JoWVVFYHxI1q9pFalde9F
XowY/ucvJBhbS+JOnedVLTULhBc5sMp/gkC+d/GL+ZZY2tGCaQ1ZyrqJzDpDINWIbSYFsLXBlYfZ
O4iA9q6fs4LA/w9UZiXrD9Tuut+t4LiYymfpTzlpr5awX3G2r6QdS4FQSqrtt05/sLyFHxmLFjPd
+cglkr5VV9rXyFZaDbifxd/et9P9KM6f5phqKykl3co5EPCcbIJeAfYF1iieu6ShtUMqGJWWpfe/
rq9I7J3G7ENxGBRNZSlzbiaipt76kFxVA8j3NH5FRB93bIMmPRBz305toljeHEzBAyri6+xWmLDE
bTYYTZHcC0+X9SVlmUmMjvBuVFOLtXyaN+rpz/hIqJ/Se7U/yoMMG2ThOQDosCV86Xe168tZ5RO/
dN5UHRNO/g5vmBUtWr08b6Nt4FpcxGmLbTybQtCRk/SSCOeQSRtxIV0PDzdtJ0VvcIKMwycMrepz
HDfeiRD+TQHP5En200xa+XqP/+uKec3QXnlpSjMmKcByvw7jS7MJjv77p5tx/yW61CgLJ04gk5kS
zZdDOLg95DL9z9sn54V3UGfiwDzNXyy8hPn6c2ifv7DGSO/oRal7WS4T4TqUEFiJ/RXcyb4yc5s0
2OL/j2/SSTsHG+M244A1/0eaK6z/V2oaCBq4RpoMZkUtQCR9oHkg+L0I8POv/iBtUERUNpG1ZFhC
jmht7V+dSOReTeaSuwOd4DbD9jWeQ3qsBZXstRVOiS6xJtbEKEiAnpoFy/GQ3MM1yJ/KA2yanNIR
dmHtLxoMmO94+rwwl4oS+3XrJAFBrGmM0HoZnMUZbGColRTCOjgRmxpt1Kxmv6yRYGXIHdjxYXCM
Kh8rZ7y3b2mNYAHAUl1NsizNXQpu15s01mzqNd+Ea1w3RfTk1deriGnxvBqwsEwNzxgZ9fjaNMJN
Jxircfc2cX4jMiGb3hjvMtEF2yT8lezu5QJePPNT8/6KmVzkFnGidgp21pclj34Rd2xn+DRun6xi
gKaq6Aq006RIByqIOmjR6pDkdZNIxh5hT1M04FzVF59Kk9V+zrKeJOnXq63cWIuTuu4TOP+mhfDr
foWQt+44hKgXE+v3ApqSk4sK64qqz+H3AVb9GG/ZPTjvUn/dbORLjwPkFZumK84SI5tMfA1LYPR6
539nmkZ82BDSOIjZ81W5HW5ccSCGHt08NwdBygviaOwBF0xHusIrzNjKmvvw5KtfsI7YHGUVfJGz
RnV4V+Be7XPz4TiYOdYCKuI/fYxTn/t4+MQIiW/T462O54++aCbJUCxXks9DAYHYJlY91SHT2VmF
bSASNIgIpqzL7wpfKkokrbyq3oxUSb+1l2l7p2GRDtBp3uuqQlfGoG1z4oK6kSFs3CtlfulmpvI6
iMWugI69j/O9qX2HRM8IKz2SeF10jvXpK3WSAqjCJaKMXZ1Yv9xnYPCucmEinSBgLCfJ5Ug9Z8AS
e+Gw59SfrDpTefJuDABMURph8dmR1NR4bVWenRvVmBUArSkwbfTiK4iLTVrTeLm02mxvoFn5hec8
yWEIbed76CR4qohDoxdLcK8u4icSI+Xn/zqpwcCIxAPmUKOZBy3+Fm+yAchVxG1Ryg6Q7l3H0iKs
PIMPdTBfrSvPU2SDmDtVWeHh/bC613caReOrxtWyP/MSpGb88exSefuy27VzILLa3pJ6pVwBGxG+
Dfs9FKFfvWKaPxBglOgo70/4ZWL5FH/w/8oyJ/HW1WR9tl58m9jBahvT+rVZV/+/S6B4jDHlt0Cg
+IZA63SsByL3FSA2TKmVVzhd4wJoMMg413h3ZNxp91W6ZreBYyxtG+7Dq9SL902IaRc9HypmWAVE
ScndTSvTvYmz2XwbKpnqk/gKQ288U1Uaji2SW/VYsd7FWBi7WKaT8TJ1+gMjR/XBKjA2hVnudtWY
+bzp04Axh4DjMFnD7vFUKoO6oFPaOsy0f/MxwTa1R/5kfMLqOJ7/lKRch6DZROXM2DjTaE5BS/au
F10y8d4/4cYIQna9GbTpqAU9TOkU2XW6V86pltuN7Rfmc6QTjxf1zrRPthToERXjl79CQK2BHOIp
23ZvLAseZ4JiujIGSQNFxlHDNbT3sXzjkZKET4CDFvK/Or8jQRx7Gjo+fsGMKnR9i7mEoO1Mi48G
8ZlUG3GuscdF6lCrn5JK9kSLSt20knZqhtHX/MacwsC7wFyEhsgdeQhR1sFDmRiLJRmKBh5HmhH7
wruR+9k5NxP1kVgu3f89XPBlbXv1xYMfBTmuhYURuQbLpGv9XFWDn7ib1kI4FvJqZm/bU79PNZou
j84ymweWYULBTrv4Rv9eu3uKa8heaYNUkeec3ztiqITUrtKy4jCGxGTXQQrchJcpfbDMHBsaT+aj
ez6UtO0TQPJFja+sHczfAbkO8wnMWTGg4x+n8FmN9hlssXrOKQE45KRWkvCp+ltnq1kxA3SJvy4r
7Y8irQsbmmQCY2945RKGC6xyqIu5poBqi6B8sPA2SQeInEMAjr7BbN54npJ6YqlnEdbHmvmGdLn8
8Y7qjmrwk6pbdsJelCx3dHylqieq2Xt5lsWcgibupgKpnRUWSvQCWRqRaApu4Lr0uwNsufbeInjo
3q9LxOIelYfvw1jkTtBxE8V++igoH/WSqN8HZy9Xreqp83NpCk/eJvNl9vtG5Lor/2I3QCS5kZJ7
p9vRBOEsrXXbE4vv3qabWUMs5NUSNkqkdb1eQol8NFmbN+QJLxzP4PNjXl8ntMCGsRuaQHQ2SZxw
v1xwMk0lJtcayFCZJgY94X2hdImRp9ivxwP1BCotUhIHzz4u64cYiJrvW82GSX5MVTaSsUcxuCN+
bLQ7vxodFN8UqgH5frczV2J2pgfm2SpT1OkQ8lM5jN3WvazdQ3UHAo3bRF3cgbNxRED48boismrX
z7+udOtCs0h6HDiRBL4JbI9wb5hpjvi7YbiakRb0r5/QJy7VRLNW+Y7UmMwhEdVOmeHglI3/PHSy
c2zz+/7WaoNAXMeZ4qNzOxrhV5kcHzsd9ySpXv8ZmaZD691tdLGa54ZzpYhxXiJkkca5jXTPb2qU
OL3p0oa5jRtD4BdKKDwhj7YFgNiw7FeIUSJBqBwWkfnMeDLfAAaPX3Xp8HNdBMQf7YpNviTFyA8H
zkQ3WweRW8fZu7sVMqqoOoRLYlXGIISkqZKjfvphBOfDtKmC+JXr8Z2t04mHbs6v8oEAfqznIiXZ
xwAz7jJhd0/YssNvETgZh/kl0hYnZyqfcIsxXXqlu4cfZ9bVZfu7+Bzlg9XvnZNT+UU1cV/WnSGi
nVaqJGX0Zg+ZTbUEHH2cWInrbxuhN3u8Sbzp9DPiz8YH05gjPR1S4GtE5tfu/GXp+ZHMWUEvSMz6
K/HebNHugB34wJ1wG/Wr2+nRTD7DJvFDa5wIsIIhT2U3mVQ9wTbzrHI74u68sn45xBy8N16GBjDo
xu2sY0srXOgDv089Xq74lxkD/diZg4QSud7y0GAGBG1zyDOtisGRhb6uslIqtgQX4oNSBxwMvhwr
tNhCYxcUXYn1a22RfoNsl/SRzHKnOzd5CKWZsEGlQ46/xAy2TrjIP+pLErOXFNAiC2n57SEx9jTX
IPioJpL2rRX/YVSFVQ/VjkgPe2fV4Ltu4aU3zz8Vjm7ozNrVoEwtjYE0miZycBVLvT4fji/oR1qT
I5cxk/WHNRrIQXlN4pIH4x2uLXvBlEJNhXTb97Mjx4lAwngKQb2qFgEH3Qw14olfZyIQMNCjEkBv
INevggXDpWCiBCDdGsOzI/EaWB4jeuu+6+BWvxot0fxwsdxYQHUb8Azjh1b9juq4mFmqT2YusHBo
f8rorJdHyXJf9mYJMLx+UcDjXW8kSgYj2jALoOlhIvrE55bqozkOwkw1pXBG7c+878RxF2ZpsGOc
OZK866pOONqxUm1f++hUfxw6SMi3tO1m4i8SucFLvK1uNOr87O4h7JuMkghEMOaQV0hX5nbL2M6S
PqrcAnk43Fa+Q0EEtHo0mmNuGxo7uoIwJ853H/VxkUgSUPvTpwCvvmte/tW+O5atJjK/JPGK1kQg
r+sxzGjOj6mRRVQWkTUerbUXpdufV5bxHIJeeAlooIInViLvO5I8fjvk9Xjf163DULLwL3OojV2o
XyRZWYVmT6HZv2IBIuQRZCN5ihwQhe62idm2P6gu0nslMpIz8CTX8+qfPnVkAOJh1mF+FXZ+s+DT
yFrGofddfssETT6/qZfsn2HZSMYEFS8IfCqHLXYdjum6IfRv8eAZX0rp6mnxI0C6ZxCJw1rFVrS+
9QW2ab+V6ccHPwKLqHv2mL+8J04AaAjntLrGHxmu9UiMl0lHuErGItj6/hQLzCnE5hC7VQiQ1Dnq
u/kXDBy82g6DlvWU9M0jpqOROKn6iVATFnlkfVLaCWJ8OHSMalcYXTOhwqc6LqtLnlcUBEwanjYx
IInyxtLM3oT+CaF/5CTVRqzxaWAQLUjs9mbm/tNIxPrWg3j71xkV+4WCv4hs0QkYIyno3mlCUnWP
IlihpHSqrVozc3DtGUBtm7h5NNGbOvMiy29EYlElofyNE1QSY+XbFlKu0fLnjU6Sh2wvlMwYoxJr
acNMMEYQIIJW5VeBNQ+6pYPg1B191BymUjig06On8OJ/fYP/tv2Nz3ERU/X17DwO2vRiPRn0UXAI
+q17vvdQhusYhsEXrhoBQ8zMcK/HafOxK6A+jpubD3hPFlu3q9WwQE/Mar6dPFid/Q6TBvBb2dqM
PB8JME4EAzkXtLov50Pu8LUECwGc104xiCeZxbacqhRKEJ9UYJGP13qMKldLxJRAnJo8IKR92LPI
O9S1CLVyrxPGVBtOgWPz6JvU2KmWmZw1xkpA6AOutQJIccyNlpCui2C1BHZOOcYnl0UfPpRgcPnv
uOTocMqxBdXGDfQ8NsXtJFoS+86QZHErqdZx+dhgVRCzqsvLP+osi5N88K1Gw53bLbHBrQ7C8smD
f/uenzHMChjkBq+lIYTCRs8+CTVRoAuQVdyKHkVzbD4cOk+PQzF/IuYqbbh42vF2/LXySK5jYsuI
S8fiL3wuOQzA5aym2rcgpO9+9WqKUemaMRdzc88/lwOltO9let2dOKBdWeKaPPYVn9725FWnaaxe
6O34prm7TznUYliOfrym/qsTUSje5uuC955z88Fw8nv/fkYq7oogfvRm6szvguR6be86oRwKf97w
pkGiD1CPXVIg9wwfOtMT9IffqRDPUeY1GQFHKzCA6pHd0GoDkjCs1XfkGf7eL9EYFn93mEjj6tCS
6G65YqJ5xfMduQNd+TCbEyXsZB5HawI/LDcfu7lDQqxmKl+Ochx6e7G8soRl+k/hDxKDBaOb1FMX
4iX1Kwj6YNYWwVVMuWE/YJx9mIk4l+wLV2foBpBvEN9/TDiXYjbRp8yGfVy7WWrUzj69BpXWqQLO
uvh4XKWtQUQFOGqp801+m6MVVY3bMXEnpWDTWCcy3V3hvEQJ6dqG1bFMSe2fJRGwajhTXI0Zj9IM
yUZZovc4k/MwDSSrDedSo/3Jn51N6T63eqil05twSEDNX71NIPCDDg+Ls1YvfGYZu0/4fFAj3Vx+
htqYo7yZwsk9VVMiPz4eLCfbG1yEu+R/V5BAK78AvYh74l3ktTs73wQRCkV6i9DzWk0hOiAsxC/x
ZUJU4/ARsZA9W0b/hdU06gufUhOpLnKXslM7Rta0mJDvCfAjaeeLKc+/dJsCG1hMjBWbK/S/ro/Y
brYjAYUXnOegCUvQzLq+TnJFcXf+6Lqk4gTXo1EbiT6qRQhkcjtMy/TVOP+9Z5epkKUeL0kuEnaj
4S64smMtsljeGPmWGEd9Eg1QptuJiAVoeXLlC6OOocESWPwLjqy9Ge5w844for6aNdFIhD7AMMBa
/IOjOUnn3nywcmLAewGBj0lxwvyPP+iZ0o/QUptoclIFL5Ks0Ki8Hi5rB3G8j8iuhRwscghMvoeI
F2+gwrOTwCGsIVBzPZqIy0rnjjSNJh1LdzW+LdVNt5DGf2MNT7SE5ogHAlYKnO7KQTURbqDIV0Gl
htsjhdstjbMSiZ1WAoD1z2ts11pethvlfNJ4YpVKEc2NAZJ1dUpY5b06w9OtwGXMp/MpUCoXz3Lg
T2LwDOx1WCO+kgJYkWioisC9YXL3WA/Wi34V5TPpdvcgB5+LtU3vubxxcIFv2R7ekvLtoUJRB8m1
yAGW4s5SHpD9lja53RcOuB78IU7oUbFZVmUhz6jZR/Jw4hi58uXCea4k3V82H5O6JxbMuj39z9o8
fjIuYwDeVor2yjm94uu0+4K82krBt3feBmNx8/R98YwJQtqM9y/OYYS7znE/cJ4/j1SEpHep5bYS
ajWf3QHLrnXXRSjM4cqyb18KOuJq5wDwWI35/KdMFW3YxXIgoAHJxk35vZsAxeYBZ/ckHEJ/SsmK
gDVW0qGJJqqQ9NpylYlsQgEBPn93mh0D6UYBuyFEoa1yHjnO8hkPDd002JVCJ8hwPROa099aB7Hd
5x9XBNLGfUNEfCR5sPuW+lSMUTCGOaDSiG1v7M7/fSuUruwk+KcdqgQklZgNey3pvpqqQIE2IRJn
7zpRwK5kRfEBUKrk/HXXWaLcUIQVRp9JwgNiiLQ3SfZ7ou5DWOJLbvF0+LCsai9u2hogBVqEB04r
rqfOGstH3q0Y3wKsHzh2dWGBRPe+1Np0ngr+7GOzOtAj9SLezh4+BbT+ayq07rUmAzuW7WBZnW+2
a0VSeb/8Z0kexK880a/itBVlgO8bWhi29FmprJVuDdQ2KRXEm0SLmYZW4s16czjeQIZzrMdzRyac
5egNcv/+wT0dMQM5DiCAjKX/enc8n34X/VLdjjkRsg2S9qmxqI5Zpp4x+AatF1aKE19YjA4/2ZTQ
pZsjRSacjEhx3V6p4DR4PcOGLr7ooSRJXitPr2TbuTQtpjgsZrUTeuXLD5cTzM4szxjpLmTa7b/4
T1oExNVx52FyleuYtpEK9Y8ds84pV4UwetSu7j3NowVK4RGOD0WDSIvLjFjKaKReuEpI69VVvflK
RHKT/f/WKA9RBK0aboTLGHmgQ1MoLQbfaGpqc9OtwESkZZKi4BO/ddZq6uZwRkvDU0o5w/LBsv5U
aLEtpM8iZ6pB5rd51torxW7qSwJ3N8SJyLICEE98A+SCDb7kgojZ+NDW/EJ8e3LjTOmLeg+u74w0
6TLv6bqqUiMfm2SjzK3NV6ClOOyKpIeGcYBjQ6mZFsUK96STHxbIwpHTwoaXcmpEhJ3FZz+/INNW
xz/XO3YK8R1wexJxmyxg1s4i+HSR4DcZRX6lY1E0Ngl+r62RfIdtANRIKDd2on4WnGtGM20SKGQg
Kc3o4VgIGE1HlTjhe/gYVny7pfPMjwC9yBuukcgErMyLDOB/QcanF//LFXC23yuHOtrVnVu0fApb
pv7f9tnT98gmUk7wtS4SwG7NttqqaZG/NJv7d7ltf6gATRTQHxE/KLBoUl00vexmgr4JsrN3wGTb
Bfjd4Irl4UwznRhiGqoq5DZCFoklE6BPw/s30ecQIwMfOYFEKqNA+NfZtS9iQZC/FKC1JnZcorqF
6x0yAm03LImsE5CbFZLOIJ8er67DR1hhjOgpQWnS1YhMr4FMNfMRArpAFPybqzd6nGPFlRe02cf6
MLpXgQRDWGVd5ia5VTFh2/VjLIYfCds9pHFE7+YZ0XC/fQ90xVZZ5f5igtbkW1SUB/IwN/e2gelN
EYPBYaZM+1BuMDLe32wRWuwfhuiYzeP9kHIzHy4pWGCPeUE+8ieiVDEUxeyF8OJlAm3+c2luth8j
0O4dSkQhnYYVxJwsk4qYCHHEg4IIPneJOIktWcpcl3EQ3A+gwbZjm9Qd0AjvInGQYNtJS4deVcKo
qyHyGBKr/tDEZ5vFfolkmAOiG0hDUVyahKAHqCAHHx6EgO2Egq1789l04NvjQMj3q5O3MoLXJMcA
jijHQeehTKw5acAbRBg+EnO4UPcskgSkkdqLpmEhH/w8v8xk95Wb6ZiY9iqlVQGsJXadFPKZ1bbB
CHM54DP9dCQP82WYMIa5G9SyOfAFC3vfEL1M84Nfpf/sK3/nXQsf/YVxIBSyq8P152zBF+sQQWxM
mhVdMg9UtChRNdMlTJkgQaJSZLNxYtn15ymUHvTmjmfYgCYM7asWYyGb6JSdPE+Aq44p/4kNjqab
c97bvbtEKTZ1rjd86wiS8QVvfkBbhK5wZ9JSF3TVHrXLJyuytXmW8svENdBr7DE8G/dvS7JYpsUW
Uf/tx4diCGNhWGC6+oCU5wANe4TsJXUnj2ZWM0zJMwnv8I8P2rHaeOt8GbCtwDDP69FyIT+xLVS2
d2RoPFgrv42SOapMNtKtVw6fFhLxOqCuRjfJlrt5vwza7XMmzu0e0M7FcaPpJQkGcAQtrw7mnTat
4YHOxmLev0T3302KTflDWmhgt3toe9BHqaFj+0q1WtxsCqpy+m3ME9zdISvjYJAR3QhhiAwKCviO
Tv/syIC0R+QBHQP+RC50VG7wpDWAsbhgxCsprjNE7Qn8rKIFwOdO9O1+hLDwHDHqJnp7l76v0D1P
8KNLRETbPoQTAHB4qVPYuB0cWqHDbKCj5SxIGWlC33PNxl4Mzf4xERiZ1VM9hdEV5aXKwQpuvU7P
dzfQWOUh1o3Qxo9SbiwPh47Phq5y8s9IzxBh+edyxdxAZk5QXlVg65P9x6tlJEu2F7wNIIxrGIVa
Bln7kAN59k+INusNecT//cr+WbIh+Ne2YzaegdhUeVFhwFCWVm41NlIL3Zao0nxO+9o7EHEhvvEC
GvJLA7eBlMXpIn3pgkVf2botHMPsEAs/QOkh3kyhDsq1pQCXnN3dHR6SUDculrOA0RuJJTV5yIQf
eK5eEoVWeQx0NczlpBt2FVmy+YUiwhxre9BssLaqQQKK4bVRBM3v0zwO95JJVnflZlK0T6W0852F
JBzWY72SpYvCeJ3XU0x24r3Q43f+OcuZ6UlNKGO36iNUKuZlxCbCtc/24nzfRm/trw4TBlPo1aJ5
qYkSrEuf7MACUmSI2MZG55XBqRqQztGDHkUcBxqkTb97ldYjW+qR3QyllmHIMGwroEOjeoKFWo+A
O0vVSi+EzcoyL+FIXRobJXkfYFNbMSXPgnzdJrKt/K8nshiWAeC6ndl5Zur305Rx7Rkep95Loc2B
a5wr8JLnCt+5MfOLnR1E6CKAQ0CSUbWA6P6zxs9u32+L4TCRkbeu5c8OpzCdZlo0HvAxu4K/uBIU
ACSActrNB0vu2/R+507lnUH6W9yWo3i1tUoyA8mr5QWfGra66B+uM7rXlCeRFZcpHtfVitKk9Dab
QkGoNu5j7JKjrKFp85FobArpr/pwR+JPHu+hHUG4SVEUxR0Ye2tB1ADORiVvQMgRacFlwbPujHn7
lmyK5af50YTWFmGPEuuOHAEIg+L300K1BvzYQ05ImsRvu8N0JFceR9TVLNMzGUCCEBVCmQeByvrv
yRSVLRwEKJfLwiduNVjXr23Gl4fOLvVG4F9d3E10o4vIzxLhojaaMBatBSIHLI0XZRaWXe+fueuy
yBg1J5MLkKBioVK7m3sk1PopbeAyYRNfUWM50KHqGlIWWe2e+ne0Jy4Aw4md4WWsCZIu4ToI/RQN
vOZVEhFKc3dhNgg40XR/wqth0fiVTjc6VOzlb/P9goC1oSJn4iSWFyZyWNZOpUh1IMQe76U2tIy2
mQOHnF6kMoQyCJ/KEQnn/Ko0ePyiPmks4kWb0qqaCCR1X/pQxKTcvjsiEXj4u3XIE8V72orkSw45
CXQGa6GGAK9fo6fZCBgfz8a2YiFA51soydIvJmckvnceZZYvPOhde3000Cs0V/4lFt2ajOe9BoXj
FEKCbsUkSz0JPt+aRLuB3FlFimLGouQflJto4ygyTTn7ei+aQRK6wfzThkcFzekp06HYWhVTFEbu
gw1ZgGaUIePV09InKz6pb3HndvY0gVXt5d+NU8pj6oVBrrdwpP5SA2x/Sr64zggfdhL+8TobrQwg
VwJbV8oGaEXWixJn0xiF1zx9LFxPl6eI6UIlIdAqYQqimBwYYxOdDABPIqo9OaY/A+kJmMXTj6BU
E5g8OlpOmT0QLBT3T9HdJ5cSGMG9jmY14MU8UOha1uwPcxR/q1aBKJ1pf22heLSFlSK6L0+7PK0R
W7NwPeUtv7RFX1jtNyrlG/gDfzSNSXI41Bdga2pc9AZz7jS4MscvqS0hzU7Az2rooENKLf5aMhrT
hoT7zseBWMaHuAIP25/exFkHdmrCEbOiP9WO4SrdZOX+yhi7LQGcEJLgLX6DPucUtPxTYGWYOjGO
GQW34Ox0kSm0eESYXhJOBjSeHSN7qdHQ9mdjscLokJIqn9jbHYBp+MGtJId2Em9Yke6FIDPbW6u2
or6Uh80EU8KTKHJcN3QTPZMVMQBK7SFZEpxSmkwPbNsmgDOmrG7QLCJIceiWxMVbA61Ett+mVYW/
82hki45n26wT1a2Y1HyC/FIk7MAzSaeRdmYabHOUjMhUN+Y5I2v0cCFDArGeGmwfB+N59+OGDxT1
7wcf5yHhWMRlmT7B7iHmoh4nMbyATqUk/S2QiJ5KncKZpKw87PIdEhpLZoXqzHgk/LYjr+1MJ+GN
08C6lgKLFt1wVP9847X3YCiDjFykvgemCe8t/HneOtYe0P1+bPyaugJ9XCa7x/GjDX341QEEJGp6
6njYjK2cbgQJNDA2HrffLd1GJswp0NMBQeqYinxK0HUemmPHZSPnajfcavTsF81zSVdtixinXn3s
x+BNchvCApOEe3XbefwZj9N3rFQaXn7aDhT6b8hTuqiJc/YZcDLr2DBmnbCOBYhlndl52d3fLJYU
aUP2EG18eBSwbnLvKwsmmotB4r439258M7sqjo3ZPVFa/Zr3CwWjk+M6Qb8mU/VychiNAiJ2KkJF
1BJkGJp6RM6TX0pkgbjgApceW8Ot0q5FAGYk35pZQ6w24ADDIomUPp8rGvlCLBAffEazqyySSIK+
GAfvyTu+3+p2SsgqQdBBjEKAIuL1tJdk16JE8iXdHVgObqAtlRc4ubCh/ArcfPIm8ucsRvp/IOgX
vMThe9mgNBRalapD9J+uLMPjdkbK8dphFZ/V/+EwV9G2Dq9X2aCoBAUcQPcHlpnogguYGyYIABuS
G46n2WKoEWi9/36ebkmbyOS8lG0SvlWM4+qz+hPwnhx0Cd1+92H4+N9ohXXC9IdHounmtTPxvc3I
mk3Un3NLhRUPC7JJvmJxcUbee2/CRn+HqwAtRNdoM8F3oKVwC9P+LKaJUKepsEYMCQhivqdUf55E
IuWc47fI8WFaLG5A6zJBC1H9Tpyh5fe5LqURM8cXkfEHCb4/bvpa3SldpnvxfsGQhsHIMjPFopE8
AepgRY3obiUaWOQkVFfdOAyDHpI1TECaBrCxjh6uw4pRMpiRsaXycs/T6oiKoRxqbkjf6nDSt1Yv
OYx4KIc1MeQczEg4oe1HuQO7NXrHln+HQLKSZWcjZT0wRpEZsvsJb0MTshLvVqpi5NJ9BbiTdfzJ
g1i309eOrFu18uPwwoANS5D0bGMKT0DaKAAZhLOD/d5VdjWIQs1w53CdfqouVvBsejOORIVtylZC
eWXKXLrtpeXmOTLpgWXueWITPyNZ8uQgc+8wUFPQ0Q5I8eFod9VcZn+Tgag8xr3hti1ukKFngVEc
//eZoto8wBJMD2yED1oH8tFZFe6LmgOfimrE1ZKc/ytITLSXOjahM/pM83q3KUop1m4EdyTTNyum
wp93vNvcItmfdaaWuKIekpVd/3LEIq6GVMf3ZrVM9IqGTAOTjzv1KGyJhsIlkha0wMwAzOPx7yBc
H5C8L1V099c8OJVX8X40rrOJPkhl+Omxi4FNd39wrs0cotymZC82x/c1MVfi+DPoa0ry5uJ2i6oK
F1P7zeAI+krhPqd5zwwKWFmGiiKLAQ+snVodCmZIBqqgKZ5XxffQd2XrpPUSPofa7XChuS8ZT5SP
iOei75IlM4bSNsK5sYiwe5+4bX8kbwI+tylBLzGXn4LqpCTXu5ad1DUabUs9ePb7VKH2ryD5h/38
IfkJOcP/ZBQjOU+yEnsbT+y7z0bhZEH1U5zq7rgvH/IsYXFUEmC8yJNwbY01otkxDEc0TlvB+bw/
qAxgR6cvxZckIw+DwNppjn0Wm9IUyLHv1jNn0sRwbgabeaQb/vJ4A99itPtktFdCPnwAVy8SDR7X
PIfNf7MSDuSAn4a4djg97oWUjvdFPUJp1sm05BCBzx9B1Oskhm/vh95pwLJIw4mYPWNy6Bc1AGXz
gkZC4+AzhaYkyywvlHEHBlIF84oLn3f3slhTJi8MTvpFM1C8JtRLIGwWqGHdlCxb1mudjma8yAPj
K+2dGIKFYtsqk1VDr8Uly5aagybl966Wmrh2WQjIaWzMiWDsjkaq/X8c0QXtEmqeKSI3eRNf7Fbi
d3fM55DAotZefFfiwdfvsfKcowcYgq76wUdt1ZUY0v67eMg52BIgGTllKFGp54+0mpOeBc3YdrzP
JqXmaHQNCUadBbEOr1eaa6YrK4ascZTlTS/dOgmt0suJbkPvhcZANjyzQJHliUWWUqPl6NvoH8s7
JtHrIQHpAeRLb8aXJgU4Iw9WMqGGLkPhPgs6H2b+X4UqRK02Fhpuo9PRfL87GyWTHxCrlC0ZMW+m
dtwXRjH0iYoMo6p3BvixLpCXVeVwdPtV41ZWGtaVW8EYEVIrtE/uS+YYDlKFMEr1Thz0y7aFqq9j
WsdzP9vtdJNM3FYka5HEsrx2w6ydZiKVWlwwoJBAaHh8dUd483BkHRqliIvTg1zgtDTgZ3cjDzYD
Ex2H+Pglr1xRGjq+pM7tof8fm+ttVYnV0gxT30yDCr/GJUL9ZpC8kaD+ouiMoS2jQpvl7ol3hHW7
iBpOnuKtAPqrqZQLtYvYt5y1urFrvPq7Y/jgBYwyEBrWUeI38MIrvobT6g7vL4BSJM2abBtDb+C9
dRJ5VP2g2zS5Y1m3MXQKzH1pqkkeRBvXt0UUI8KvNabiPX1EIpfe+fpW8CkGPFCvt1JmnzcmVssH
s1KZDS65bkxBJgMKY4XLJx8q4Oi8uAnZCWsiS/nx8xo+nVRM042V+saIEFNzgX4NeB0CIp8r2+po
rd0T5r7U2+zk0dp+qRj4DEkO0BjbNwTFeaFZ7HPFqeD1R058a80rUOkWWrFhEEcdKNBWmOPvc3Tx
juSdCbdM+rrJjkV9sRbBYpym6EHiibcs/o0jB6oiMK2Pj0QzPZSDNSsHXTQK+W02yacctKqq1ceW
fhDr3YYnibVJBSmkK29hB17boOT3oCiHgn2MqbR6t0nkUMP3HWcMm4qgYjiB1c91IJ9/4hzQWDFX
c+r15JfdX8/NfWvz5UFdXKAQLS/xoB1GilwJh+c0QDBjjqTE+IZDXIQwfcP/riNL6sRGH8bdI2hR
9Os3aT3/4asGAw28SExtWgwDYVkbcmuPDtBMXvJob5DV2npNar9Uj2OklRY9yUnlUwPboJ03qjwI
2aoGj0h+CrFgwsLNRrQg99Nf+cmPUM32AzIQwP3ufRqJ6T3YFNQYAEX7OkpAr4b5B4M8fav5Aewb
QHdSY3id8d+aMKTE5Hlzgomc6MjZgbVHnQoed2zciDaODvF5olx4YYgmCVWzbsyO+xkbPqobGs0r
KViz8sD5C8X9KvkkZvxOEnrGQEuExOiaEFgP6BuQcJ8NpgXIZC4RivkK4DsCihwg0IH+ALt/qtCz
P7F1KbEJYedQ/ZJUpAN+/Mv5RsFEhLZ2u3pAyahu68SMR2JxrEXPeeaFsWEP5kTtZHScs5qT+XgQ
nTAaRctYiWoGvIDsAfcw9iLZJ2LYIzpBiyNgKw+rCfeFMDN9SQP0EEoez8VQ91yei149eQnT5fpU
CUIIK4tfA3sWPlqRc9r9nCF13ixBVOW7nQs8ZJu1fTtx3Abp5h1ZqsOpzInYL4su98lguyOI9t2E
fKZNGMj+1EcsZ+UUUKmud/hS9JeCuEla0cmFjimMFjWktQ4nXo8PxnzUlgVo5HWBhXtCrpKGAh44
TpdwCsSsOxeKjsgjjqssg7HJNWPbE/U9LNhNE92RDrdZtPEFGQPrDYez89AuEjR9kLyx7ElmCMbD
fVQv4pa0G4vlNE31tPx960M33GsTSsl8z4fGtbMRT4h7MO8fg7hRI/0uP/F1JiAeKKhNAMWUJS30
jNFVZKppau0FqbkJ8hfek61SR2ObbPJ3YzVNXs16ebiv2tmeo7CGflVIJN3THJEHONqRA+OV3bj2
lS31tzd9F29PuDKuruqhFBkDHY/tEfWWorz7aUMX0rep+eSgA8oTlfVluJwqGNdiFLkmX1GVONwz
TKokKSWlsOytfP0bgsqTpyxSH+/Pkywzw+cGCQbNoQ5/OYImPkSMKPTyLUFnsRqlLldPQkZWXdJa
8yBegrHE158DZzvh8MTcavCZvXirvscNnEzqfpclQOWx9GwEMysDTQipDR8kc0MhLDIyzQu1eAk0
gXQtv4kL5Z9VrlKDCeBkKy2n9bi6FSkrhz1z0+C43wjdiH1o0KjlQxkW8lyjP17kXOJQa7DxcNDo
tM8jgVCdWsFSkvVCviUBSyqAV7TVv0qNXXT9gbv14jy7PLqlgUBiZKt3w3/ARVz5x06AkKnSJi4P
OEDhPYnNMoSLhL0o+K8bNA8+xfMUEUEJmxfI08OIKzHw5P9cd58rjV3b59tMjRI7XD4KPZiWtXAE
Mv/BXXg+Y2qITuZu6QwFa+YmTN0wlkI8Oit7zHeg32vpV+SYJSvZdFZgnlWXGbOwfO/o/qTjBmhW
Oi08fXbe7vYPKRUZD8KtNOEUZNGSPaqJY5+lBACASjAcuRx88mPbaKNypt2zcZrFdsaluXPCd+c9
qfVTVDG6AkODih1X5JYDsbZKCucE42jBmJwA8qjdPrgCsC68CdgCBmD6nUU2EL2PCC5fJUfOny85
G8nXeydM/5uoVEogaQwLjXg2YDLhVMXeCTjYaa7IdOVf4KecntZR4eGM5HeGqK7doJ7MeaJOv5Ha
2IVsZ6mD+g6gqFWGxJgIceMurmZs8JpoDzHp+KLYxPb5JiVycUrzztQnD0TeamhGKOyogXmFIANe
g1M27Vp3JP5BAgUfJcXTxrah/Fl9KFgcfx+2hmA58BpUj7XSHlwoAmBg23UAW1aHiUg76JLCBOF+
MoDlXxvafcxNAZKhSoN6MsIDEdmyPj3zNw1iEuWln+JZ/8kTnTQhv1uQ9vsORhmiV6+H1ou5s3xL
9P9NKh3Bb7g0jf9VQR+0rbwqfTDbaiqa/M3xl72WVLMmjfuuHe1e0kyhRFjRKGSnYEZPG1wSBWuW
ioMzs/vtCe8TxtAWPiYqnxWNmVL7Dm1cZmjotcxXMSfGC9L+GhIFczCkxwRBcN6Pz/rWsumjzLC1
LOpo+C/L35REyyWi/BXjdzeC6lF4ofAfEoI47voGhQCIWOlRKEiGG06eYdxsSmac6RRlU1C7vG3F
TP2JqJNXdR+qXlP6kdoKNV7FiKzLTMIV5z6KM0NQ6DWJMppzQbrMfbn7ZDMV0PYMvsM1gSJoORii
A98uweyrazTEwtwDeti0zVuZY280Zy6hXZU9NmSVt/ergfj1+gTc2MtEiAhB1d6hXmlL2AfjD8O7
eDbDaWqMxgCdxNXohLypeeDDd9AOEG0RKuL8pm6d8FGBE2F/nioyFqJ/jRDFhN6dXfJ/sNkzuC44
9SaNtGWUp1oCMRmsNEe7J4XSyZUI/cdSF6Upzg5cSAffNx12zf4qfX1RWGd7lr8vOuT/CfDzUIJi
iMlYdJg5aI4vHj670FxtZdH8pJR+CYq6GoXznDhmZ8wbiPlkyY1Nr6TskZv1CPQeM0hgWgZSTGW1
FijdK2TMEtf1s98GJTR5CQhArsG1E9WDRAi1pZtzG7qgmaTmaJ/MCWmI6QdcMG9Kdv9Ocb2EgPqz
nfNpJ7eXiD+ecZy6nwEjIP+HzvXJ2n3bywC54YPDbqoYsIPi5kNvqt6wmgFhc5IzJ9suL26BILEY
f/I2TqiHB0Vx7kj8NXH1fT1k+YHWXJBUvXE7Y1k5oYeE+2uG2QIdugHvNXbhn7ktbCmjwx6ubGmK
BdHwyzWSqYAYDynzt34oF05RHBz3FaMZNfC+zSOYBt59fMUmEEKv9HBBb362PC7zuchIw+o3NoUH
QEDgCXYjSBg0tHDrD6UMoIPVwvLQ0tFwlDOGWq4rYXYGtWbuOGy4NTq6OQg8BW2iJpHQYmyP+YfX
QCUMX89k/sE/ptPVREd1mL6i+qzk3Fwh9YfFE1ZckS+pI+k+eUhn6qXDRA2klpusaQBIDXZtSbRP
dcTgTbaX6QLTbQpu3dUGk0JDcUhouTcZrHTRiatV4sGPUbAfsWqFb72tLCmPlKOiuQcneJuGmNk0
6UpJzYQlUvUy3U6i7tsPfcFnl9uRL1OuyoXmX5OGIoTenOFUmFxIHox3oX1kNctSnTGm8gqBT4CG
RrsWhXvvUapbdxYZwTdMHxtOSSy9hfNFGcqkjCnxkSNT/D9n4qbCbVut8gpWt7P916dzrB12yFC0
kAtIvda7wWwl46mdao7A0mopFQQr641ENkZ4PbwM6/evOk94WkiBtoJJo12uBBT+0UAYx3QfrbAV
pxP3521gIg+FZXGLTwJ0amcPUZ7BnEySmBQGLzAiOEqWYPnuIEwsLcikwHu++99/KMVZ1pmdx2A0
kVO+xDh0D9GfuN/PIUlcedg1bs3WkXTSqJFbe06bwyipWlnGYWml8uMqY5XLT/R2Q0nApDm0VhfO
f14NJkq08LWxFAblEM0Px9KVhMwbyVutuW+NeZa3l/vLFVvtijt7JjGptCmqrtPhJQBss6ivYUAn
bYQj+XR05+4O154+ExR3PxW5dkwJjpalBKpsec0SMBN5We6QRCDtn1mBtCGT/hTGk3QejOAS2kpb
gswzdfdMe9hfVX2vYt1/5CKf3MaW1i5SkFBcKmHs4PzuE1ktXoc6rBhavVi9wglJTegvW+SK/9gU
DfD6VHjBAMpXwyP0Cgm9/6gmgrmOlivfm5PmFAywXjzJZCh7cYRx0xso2qRQAwqZmoukGRGhKZ4j
BFOxcJNbaPE4Tr9r7pzOGekZ9I2gZiCOsnkDML+sZ4R6zumNk6olKo5H62a0zGPF4znUW+oJ8L50
WF2eXby1tsyDLoYvIcAOw97DwoCHwcLAdhHpo7iD08+o72jSViRaAiCmEVr6ady0fw54Fn/aKeue
Iho0+n2Gtd2QKYDJ5RUa1LrV1qu0jiQ7mVZ3EpNfWf6dUIPXvh17gudCEQgkP8G2mYTx9ZugXM2Q
ETnt4KlIF8X13A2TMEbnbsqbHqmRsrIOyEUUDMjIACI1F1EU0A4Ocw9IB4XL8OyXTd8Rc3xyjDkB
vwuln0HE6sn11Zdy+37vljQWCHZS6TwruLfrQ+dzbU8sWhp929VNG6NkHIKaT6bZng2qrlTXCcoZ
SmdmBcE/aO6dkG1FEORERkWOiU50spVTU/QSJhxpVbkRQs8ZyW6g/gZ5qeiEDwWkIjWdq+EqX80C
eBWeWj3cnSccufuGfhNcCxeLwe2u/kULICaxCw6sVdUN1I5HIDZLBTYYcLeXcT74mzUJ8nWOkIGk
ReQgmQgq6Znh+/2kQLY9QcJEn/o5iKSicWF6mwsEL/bmYCJJkuErxcb25TR/J4Ck0AgzitoevI7w
m87c2pZBd+6q25XIT+BIet8pnxDruluZGeh8Uh12SEanpAK4Mr1EkxohKL7j6LlXup8QcEFtYop9
mn69JQj8oEKs6Lca1WLGlmbk8UNborrL+4kgcor9OcEBRXzriniaFnq5Yv1BBKzBRrAinBMNAVNY
bJrn6/tsme+3PShwF8NdejNRM2eYVR7PkviWEpXKhk6EwQCaqhBGeW9Y3m+sy4NB61pQo95ngReZ
+CqMyZ38ZayIWZLzqMuFa7AE8HCjzNwiJhl/fUacQHV6D0QLPmR/KQ1kCRISlJENS87QVRLHVkab
QK/DnUJcu1Z8eSXnapW3V/rhjkZRFird9k9UA1A77pryRrO+qTbk9r0ckkvfPApNgCBdZUyjaT5A
C/r5Vtw2WBTYFXr/8iG8xY2BW1tB4oIcJ4DTVrbrCF8mVtSVJhJ4SV9FOGSfhY4vtQw+ka7UGD7r
w8tUWvgtq4p5LQw58aLdZyr15YMthH/OVgPNlU9zSbxkW9F40Lpmk9FyxsUA7tRouJbl28G1ZXt8
X7EG4PhIHeLnQxHTvhTjTsLmCZEoa1XYwXzJWZ7J5ke6c0Q6c09H0bUeFL5CC/4igFVwA/mCRaHJ
A4X4R2T4b6Ss61JcL1LeOb6sBvQmADhxMB/b2Hm2F6VLyO/dOhkj7rgvESahAN/yAoVDp7uq3hJ6
QUhOYn6ZbhWmBMa/Gm3dA8+GSyi4tBIHfhk5W5qg2SvBpDZhhVEDS3s0WiJrdJtWrCSVHShw5JFd
5FUHTRF5dqxTB8LmMpsrdjUEoEf/erJctFkRnAE4uB9dS7qvIa58Yx3zvoJFmtTN6amPYoDF8QRk
oou0HSxhDsSokNT6hCKIYYdQI7fCgFtbHAlu747unw83TdPazj+9AZxZOcyb+Dr/lFev//qIJTCQ
9+XMgTlCTJPtshs+Y8kYdBFe1jYuGmENvocRT6E6ToQxV2R2lVKDVcxHlUWVp8fXG7xaEgvxxm9L
RiiWY8Z5cfw3MWsc6ZN2l1Z1r4QrIVuz1MWSAaVkj7vYqQ+2MvBAhBumZBm1gKsPPRQh8JcdHqZE
gR/AdXya1Thjerqzm5ELavXzN3QMmHOYYjvvRmPXFgtWapJ+O/+6w1qbVcgzjxcvUbJewgANfSLh
GLx/dIuwp3WWHNEElg1IAqYYVF5TvCqQ17xDPoHc/8ZD8tICHo2ZGVFCvDzZXPXm1W3zHAyYJhQA
OoeYRF6SCFqdkPqtOEHEQJDqDYszpmpzjYy9kON7QNzs3r/BUXWZTYxD1flOwyqdpFqfa5x8NeQi
7mdVyA1eeCk9FKkEyk76bc8Jt1uRhUjd1I6sz9Lwkp3z4YOM2kP8AyB6FCr6FZ9YNAT8o5DmhbmH
DtUODlKglIc0yhObb8kAwcKh3HuHfDgB/+QKSuuL7yVkDqCYQSbjwQcL9T25YFld3/gZcPfqKv2Q
XfczRrsQKHzM/pfI5fhCRrnfq2wwPgHShh4RO1A7lQbQTna6JAdYBJmYIUo+Fzf6jXBG8rlqJFmD
9Zke2PjBpqUcS1EEmVWs8HFdHjNgwXrs4PNNitehBPUrJgDsfweuF3PtM5g6JlEUKO5BcZnlF3hG
eFjor/r/BD4zREF1FWs7dIfsexi7b+fquDFDhkmXuP364BKEc87eQ5Cc560SnS7Gza2Nnw8f6/bg
Fs8T3Op9PADiLXc27J035mozGooDbQk/az6VZTGXNFwncUegl4+PCwdIXv6pDVc/FKzk6PEyJU4O
Ta/k6BqxTPFdhfLh7bYTfsDYZIu2X4ttoVx80pV3NtgdcH0g1adNRPLEkhNqzcfEKA9PRnD+N1kH
PNsKZi6WS8ZB/0c4U4/UwhF6vHfTPxl3kHDCB/cMq72BrBI6TTtsg/wFGRLnEDTn8bRQQ5oYzkHC
lwU5jEW7ciaE/x2s1p1mMYf5/lc7cMfSXuhlsx1b3feNqje/7FZGyJkxlxgjXkZ52S4L+1HVmNIJ
ABioQbacQw+FGe1KjYddeJBfnkZxsqH9g9MX2fMWMpwnyKhLpfJ7v1bg4N4j2DowI4m0y2dLWDDR
Ap69WKCncjQuNFSrGKSGbvwtC0UFUYYiw2d1McFspgZ8R4tCwYzHFTW+l52qyjJlzeRhbv9njElX
vPVUS53+Gslqaf9l+TEOk1RICfl1ux0if5tgzFDCDeuqmH9HdOH4oTJui32kptEUf+gBRVw+AZLC
+/FAT/DxtkuK8ILw48Hyx0fT/DzH7xL7+qRo88bfXOBcMYVungvWa8ttk/dnr/6ni9IzTapI7MXl
WHkzpIhnErD9AZfNEsYaSv9pjArUtUaLeXcKofCYvg3x+ZMZ1b01ul2LSzX9wdP5lOdO/uLMAmFw
QcAZXBklM2sHGoVRlsieywtCKWOhY8sj0XXpFnqXQ3M/N16D02pfct6emcvGI3WKCsNQG4VurN5d
RT8XDULngflwxED6ykqmAzngGEA3luMpDbha/BXao92nJHq2plzGXbfzjGGDmLVslujf4GK12WXL
7IiFYA3WTpJh7At0a5ZK/qZbI/zBoFZ/j18UOWsdxDPyFq+ExPbt61L5IJg5yjPrip5r+pADrfib
7YS1Wj0Go9GckcUNBs0n45BI83O8OPVS0i9F8Ts5JYisOwKG7C5fLTm+0Nh0iEl/xnnIqyUSbYFr
ZLpuT2P3q/3uQm1TjM3jsiSw0XTdd9CUhJnY4SxeU/o5S2WAiN/aeK2X2hUTHfhJl7fIIwtCIgmy
j3tVlkqRrJUBKPE1fTEXZ3LDXl8COeIjlV8z80BFjtg0jP+FtsOVrWB+NxiNRzjqzE8Tpu4+Br42
1JoPRsY2EQgG7iJPs6WcnDgGnn/7VjpiywEwL9AjybintHMnL1BG0n0dhDK13Pdzs9T91Yqdi0Rv
XQVVJ+zF20Dx7RM13YJRkrdA6q0dyW+OzIj2bL1n0CeKKmn4d89CvBW2ONJT2hjoWPUMB9E+mnZs
lllDRCoXknGmk8a8Z2xuQDj5ohH7xA0np46DtsKrSnw5uSzcijg1ARlntHy9UkWZFHb3pD9bwoQ9
qEoKCH1Bru5i6A9M2Q29oxLAwgoLyanBZneoEEWBFdg+9xYInPgv0Gd1rW25Aa7i4ga3SoVDynr6
eOKLP4AuM0V84QEgIfrGrT3HuJ5Mq5tIeHFu4C4RsDNrarUuXgvHhXzZ9JZidrrqyF7dIe4QVkWJ
C3FSZvV+kY+EbfgpAY1TslZElUaZghKV3o9yj5uWdF+SVS8a7Ze14oz9vjzvH7rdNIcM9XFJ/vuq
EnunMdJVG/3EzHTVyGJRM4r2BBChHd/xlZ+uYnHuErXMGqYHnpNcDBuuRGYSlm6xhF1duTR+l+Gj
vYO+Nd4DMsNSlmlTWI2hpDpEosPgu7im5DztLsiODXH97UGk77zOqOw1kq2tWPFP84b2jDTV+C6I
RqQEWl/+vHgjf9Rf+apiD4o3yAr3m1bKJRiWk3AAFzR4PX7v8TtY2EQqlog5Q+qy8VE2FTDXkAP/
ssH/0xtyk8eA1bYIEbnQAqJ74IR0sfCsUPV8mBk3KRV+hqTxBsp+8yMe50ZMItDvjehz1A+jzKC2
f/mbvr7xczWZ7JoxlY9KYe5t/fjK1JxX4tF7WS/tFPRB182o7ixxA75UgaYuEOfkmJndY2Fmdw4G
6NIg5kDLjfXNj8Rc0tvrg3odgX8MYw1MrTDK1a5xBi4gXOrC8pM45jpnAsFYYIEgcbiFvn+CMKEJ
e9rbcQxghbqlRdUvSf7U/zSTGYKPXX1mOjH3pOX6OFXowmzqMLv+188fjCjMzXZbm5ppy2rTMtBP
7Xw9YuMmhxLglbH7+x9Cp64QwTmyVDSuN0V9CxfNn4dcLOhFRD8SywKMgYZzIYZgqqKQiDeSwxM7
UV1YYydbbqUTkUM6n3nzlQw9KYT2UT47oMIpH4pZbYyUns8mPmemy9V3LgYdlgGyr50rpnXgfbew
wQG5SXqCmtBTOYmBExDmpUQ2W+ONxRLzRi4l7zC4LR5qxqR2N/b9M/gFis+lmZ2vJbU2QVWxph8F
2X23+LFOfq4aqmuYx9e2ZdflWMCqKREIiRr5SKxjJSoZPOd8G6WS6itXP0AYPqWQ1P/E59o+Am0t
W1qbOhh/p4O8H9Z36nhLgAzQKof8GExuJO6F3DnYHRPOBEivpBHfuxLmewdUohtoNzgfy03wi7uS
KC0gENbqBanmBDXnyRfhMQb36Dqp9URyvRTygD5/zYfu8WIzc/A4gM9mDohvSNygiPPOTFfebu9P
PqiO3iBSl7V3r0lyrp2VctMfeht3Gq46mZtjcMjTB3xu0dTHR7pST6jio3ed9vlxrPWMNzP9/YlM
mThoQ+fYelgm1H+3Ug16KRhhG05lvNaq1Yc2RqUuz4HeQ15lYiisq6+Xx+/12SiwMFKO/T4drH6v
tViGH+z7ikS6aJDqNzEWgiD4Y/p48i/J4D1lVsUM2+j3ZIa5YdCmZKRw733J6g0Mv73st5Z7ZEA3
6pXW/VSvsvjEey08MHLBzJYUpyy1RO6bf+cNMhYJ7IGzGMJeof5sUKjc4/S4L1waclFKm4sHbMX0
jk2o0hY1jgcqp3/vxDzTXHEwvyKcQKMKqfNvsp2XCB0IWQqGAX0pPyPci3YuJCb5YORfEgBgeZgB
jg2cxK16dCYVYjGJmgIKwzaqFiNKD2dfTAJoxoDaZh3NjHb7kHgnCaHOmiEC0gpKtv3mOpKDxCSR
TaMeG2I6vfRigyNTnRl/Wk5Feg8ADypYn6agWM0nxaw1UJGvySDVOpGuN7BMysqBiklQ976pCWln
xAqf42nNO5Dn0ojGSMUzfbjUQ82pbUxIY4CAy9flYSCV3UA426Dn3GLaR0/fyL0/1BQz5Ph9mhv5
zPc7CbXdSP3qnm3pWH3yRW9JHP+dY2Ulh6HTlDZ4FGHvF8JhGaz/O42WhNsAKZeIbUNSS8/utYul
NqGO0A/h0s80veKSVD3h2WErbUb85th7fNwUO/+0Mvuvfv+pxnQLwUyD1RsOcI8fU98+En+m7Yrs
vTh0XfIeIIHAzGDWSB0ZUNn1zQ7VbYs9YheEgfvdrQhzU3NtwUG9JT5PSilKI5Zz6df/qruIiEAB
ojPBWfYgcwlrJksolnSR3+xqY5SZhuUaWFlf/nCI4/Sroo1I33HxnDLe9nwI15uB0fCAK0eTqQ+o
IcllkgqSicRyuLYlvyqo3mP1Lj4A/bYKvtx/Cgh3GfSfqbeoCnCk9lH+G92mrOaVGhT9wKz439vm
vQr3Z6vYPC3RuxaIrI/+x7TrdbHfEY12COeHIgGGMv5LQO9/QrJRcRvTgwieyK+7oVmqN5fUKC9X
HJJO7q/GhlVLJVfzUJ4+DdRMD7atyRtOHqR93wahmo9KvUaX5Un3DFQwCn1Bupixd4ZDAnCrzZxS
ziXdMO/VzzghCJmMaEtEVdlLiZgvy13rCmkuelqxKmPwBDOt8OC93tLp6hmdT399dCZY1TQ5eIgb
VcGjp3EKF63DKwRLfn5ENKpL6w172DoLPblmXNi63Z18Io1lz8RsKVpaLjWVMY5jKorN8QnHx6oE
utD5VntHXA5TfoxmXPAKLBg+54ttivrLvRQOsffvIma2tBZamEVPPhvDhOWgMFizLKvFmlakV5lW
u/SZLt/SGqOYe6viBD4RgltPpo91m6AlLnpR2GfO5G7ZLVnmxmkn81ecf99zKXtdtOaukgI99OEX
oQG5IX7g8Mg5qGNQ4GQabZRs8A7b4536jVDjQW69CQLJnlviBJlA17N7RhDAeHG0kBiyvaKvTPpJ
JIgfd2b9VU9rXfoCbpjXCyCmO6A5g8uLQZPEkfMjXBiimxfeu0Hc2TgSqduJXjxpCpbqmZvtmqw4
nRjU9htP7HnfQoY6XLbsQTGNdrQQJn0ow9gizUXisAh8Q8nITHb8Hy4yzc5aMyMJJlSRIWIdH4K5
me7GR7lA8ghmEtunoDRpi0WYJomaNkR4rneDmn1Y+3Puh8k6/Jpy8DdvfuAVTUSzZGy5m15pOsBK
L9anPS1Xp7e+8lmBDetaZxQ3IVgGaJnI5oOMYmBk2ZJt7Ldhsas3iu2ru6ajrJOMhir2jwrTzaXV
oAL4mAQwUSUoTCtJvbI2vWiQJBFv2Thz0VMcCiTG8wsiAafZqicPLePHjGShcJUw5kgY32zkFCaO
NYVBhiEKpzQ5S47HaoluWev5il76deq6OfT5XQl29jT2/8jZC4pUtdIq22tJJG+KHjWrnpNWeAyD
4NKXUPlGtJBJpwrkk4NGRjcGHhhxdEPvhm05HXqFYdfirJuO3l/CZMRWgvfgLRFnDSb/5JYMo2lU
qJS1j5ZTvbtrA8FD/CVKtTjWVmuZiTOb3BoO+LPy2tJHccjGppziDjIU34C4kwSn3oFgLd6uwJfc
gsS9Gqi3/Mi2nShkaCSSOyXMPPuKvkCJPREmcXCFKErW2UDB0vxFH9SrbFqo9dnQHlThx64IqXov
h+FUcijpNwVXe1Sg3K4TPPzwBFfv8sP9Ps4WoWbFbUk/vYaaEho0LIprJoeBdEu6Nl3GEjoiuFh7
mCt6UTGBZ4B2J2wpRLEa8p8qrZ6XnjSwJqsUlW8FqAzbdAjVrFjp5/PPXZwcwDiYxM97DQxNsF0L
HZpD3bar7Zk1SICokeyMFWMoIpjcUzxdiaX6AhWvU38Tsg+wD6pHDT6Bs/xDKbxhGp5HDKq1jXv4
Eyi2ASqHwt0+aulNpxlDfXvJBfs1iijkEmk5SzeJuXwhDV2yRfiUbhmh5ncZwUVZduL1d4l7FTu1
tvOdlr3VGHMM1quVAV+O2pK/c2pcEtsJB5RPfghJfGkOcPywxEhxzTW6KLmyI1nnBjG66gaplo4X
4gQiq1bhIY2k2z4uwy3lWz9gIvOJMkdP0mtCYXCsOLH85YHtaepw4zLqrwe24GaoJ47HZPQlhKvS
VPI89vfcCJpMn2wtdSudTRDrY4klXB/scxY8nQJGT4UnZ+Nq5a1CzBzoRbVRBQTsuRoehyUK2JUK
Cqam7NqNXdNiclhYrN5kHGLaqoexvWJ3bX92AgmZXnQcVVgsb3+ioHaEbMvFAEm063UDogr4G2gJ
P/x/iZ/2V1+BkYOq6K8vf+pjBfXlDKRyOX/Ariq5fYQ3LyB4UOzOdXtrZ8QB2WOayGFxqr6BUV4e
l2/A6SSWh158vb+93g5iH2feLY+k7yofWHz9Gkv1jfACso7zwtbLUBH05KN2QDwYHHiAtCZixQpP
93ulFYgiUPb4YvVZBJHcncvhaoAbniktH0T5vEMLLdJYJBUQqLR+Q0L2eLulpMME0Ajp3cqT5oF5
WBbPb/3V4ef+htFO7iLNEdRVFS28A6rHC5bZKUAEDyVuYRJdCdGxY0BRh/FWTidd4XynoGHWS/G5
LzdO8M23kAt2oNTe8lOkF8CusWxxwhZt91yNWD08qfqysargYDzLgtw1sPu+/4LyCwkqFehnwu4r
FOGWY4gs2F1wbarT+xT4glEVDT+6aH3+JeRi5oUg/SfEjh3d9hxQIYX2qqKRpc4XyFzt1QQ8myi+
YXLQp0BbT9f36hHbJP9eyeziZhWpa8GD1heZJURe6cEPYZxg7VN5o1EQED1/NfGhYoh5ZJjbYQuw
nSAMs37EKCksEt3QnFMq1/yPBSNJztvLdafP0xGadGUaV+hUFG21TEZ4OAzKw1dz15XKpCXfQLNx
1laL90qyhCbSHUyOSEOcNqvecPK5SgZ6mesh6kJr8F0SQkTHdgVSVPXAbXt9F2vpBwYY14/7q5Bz
jAbCcLfM5QLnyVpy9NhWBWRzUAnGCUpjb2oDQ8mV/5/GkLN1USvhS7N/BkVxGNsRX0gIAQxNXGo9
o412rNy6cJov0GmW9CC3AkIJQL6rKle6UIuAdOoMTdVcHz2oXScRwjflwXz1Buj/d08gZlm8eoLY
YzUC5SK/MjGpa8sF/h+n+8nG8FpvIAXhuuThTESAjjv0C9497EgxU8il19sV5ohhuEoRGf9T8zkN
Mmy57SWxxHVCPi1025QkwhazqzNWSzPtEYzOES9Cf/KO/L5QtOVKd5NRSaQITPUZ0fMd+syTR8fI
pDcMCtnocourqPXunxCFoGKzx0JAo8rn57FxNuEt6tySD1KodzdKx8CM6NDrd0R+e7rvsS07UpiA
qRLRy4nEbY3YpwyKftStip3tdj0759BKCZRjQzeTRwI92fRE9i224WHl2VNjG+r3aTHi1kL52eAz
u+HVV1hSfDUK1gaZGUtEahWFyqT3L/lA4m7oEJTLMuCMwMh+O75wUizHRTcnAedO9TEvGwvbYbg/
QYDM1MS4X/Sbbx6Alxxs4otwRDncgyVgxHgpZIUi3/KQVbdHh66MYoQtt82mG/qBT+eBfGQoa45V
G4tVMPStltcOvapzhd02Ox845ptljxxxqKddaTtYKhLYJz5rA6HUaUajqRKyJo3DuM5DEOjeXsam
aJ8jDrLVzdB5ShaUU6SkVoEwdPsjvEAASMwOSXuplOhn/ZbXxhXi2aSorEknEJftZ8DEuM44caIQ
lQO1m8RQFs35jRb4lxGprCKkXt9fraTjWBbBtat3ghg1/5O7P24qWbz/AhGjWRJfqSstNuamcFKb
c6VB59H+PKErpXHsnpRWAIV8ibcRGjI3DZEhn8QOkcu0MkrCJkbMGOGEpBRorlYzFTzdiqZ6BAMK
EIZM8sHvejHGahploXdfFMw7E6ogU+vm/L+OehDcPCNSv4XEmrEBblL2O7Lrmw+Q+ojIB/4vLFL2
AM4RARKVb5A/Dth1X4Wdiq0/E7oxpT0kQHmv/yWTSmxISjKhFhlFfP/EkBtn0KaKEC1g3Y5WEdvT
Muv/75SL2m8ecuohDf4gVR3924JvEJdIQtk1Qla3IKJ4sFdbuo/ydSvpGdyWsXUlEvtM/+6p6aLI
Ilq+xAP/B1/E0KGFVtHk+WvhOSJ6vKENXXfmCqkTrA6Fl4YWvligllwWDFO99wN9IEX+uaRqU/Dl
+YZnrQ+KIEL1wiVM7hGoKRwGZNnTjDSfiVBRpa2Rngz7SnJSGEJIMT84JntW/nosiFrolq8Dlr2N
NoZJVrBX4pL972VMoL7bp5V3t0jCHZnu5WGYnTLGHrJrmeXIpsZ2bgN0PBaXQrXMdQK24s3eelhD
+35sZrRWVx++TAlz1vKrBvIvEoX4/D8SKeTAka6Fyjt30le+qtWnuwGWAhyLOerVvzB+nZUyk7sC
TywXfG/BKA43n199UBb+D4CS/oikIzMg9pYr5CK6rAfb5rxVqrqBlNDN6bWcLTPCy5nXGVsx9k31
Vk0m/NBkG4CkZS4RXUsoV0Pz13oS9KBLwgURFd8HJiuLB4E1OU6BrZqz3t/nEEN/tCjQzRDG1Biu
8x5+4xqh0rGSWSJ4sFh9PVMKn9E4BYYXWOTppfbUfPBtMMmWYbzosDzGP/DcT+PkDQa5IqopTCvt
8V6nf0sUMmnUa0KfQErFS/fpXoZX6d0yev+EKh14f/U64/G645/5VWP9Psbb825FSbcu11BBgSUs
Vuepgbi2Xonm6D2X7tRf3zhYNAGxL99aZz9hi9i/vCY5ohMaf1sNbeUOj9lEVE1RgjMJJOAI6Sgd
u9FEBL1zDnrGAqBoVbKRTbHn+M7gnM3Ye2d3StiNlNW2ZuEsu3XqG1xLJUY9tC9c0/b3Tp111wL4
9Fw2cSt1FNXL8dMJuZZcZfN3sfx2ozNxqlf8eeYua2kcqPEpw80aWHVQ6nhrL3kTL7M6TN86nXEL
PEXNX/nisOPN0dsUZHbCM9WfkwhWNNfIe0JHbbXkn14alr1HpiPaVAD2BGVg8cYv6FaBHJ2HLFsU
mEKwszwY/04GUPMc3f4VvOhA24xGv9Gwfp2d5GFz0O0CBsjnjU3eQoU07V61GA6LwPkLIfVh08Gx
RoAB3uRcT3nIsddvLmbnQUG4YgW53Wht4OQXtfnWpYMS3xDdIWQO1NkTn1bNM+7TVWNXZbKPp/va
iA0ODKkKTijbOYFffNQJjyYYU1gI4sR2p76VUNlN6SqER6GeEja3yc7OJ3io2K1M4jEcv2l6mkLs
Btg9iUb3204rnVpye3q8gFW56wpetfwQRVg4etr6TxcyGfqq5QPYrWEImyZ/eVOgTcRdJUweOICW
lNrlCDkfBUh+ORn+zGt0a7g+/tkCDfRvxLYGksAb05GEGKZZ71VO63/2+WdpWfm242a0whzSSVFX
mdUhkDyZL7pMld3BJC+tINvOKubX1UFB8u0De5TNaL9bVnbV4gKazunVGPSf4b4WtsAPsRuDVX3z
D32JAf8wzzg34C7Hp7Wtcz/ZOL0ShLhj9iVoTayE75hKBimDrp28ELsycD85/Ay+4vWobeB/a3N6
4vvA1OFkxRjZeW3GY8xA2mAZEuogQOaR3SRGM5u+KQw2CpqNg99SzNEHjeRYjFo/xDVve45s4na3
gV5z4v+Q20faCmQyDc1SHy+M7QiGKEOdb6jVcn6EA6mQnR0/5FmiSYoUfHNkWOBqwVRCuGWqIUtQ
Ldkv/m/28JcJK/4ror2Ki1kNeSGZozXi2ptW9IYm4e52Tm2kLE9N4xvLagXRuM9hNtGVgYIYw2Kz
wp/fB9XrH1/M0cUSb65hZiuwC3rU4XfSYLzjuql+d9Z7lrt21Xf7zQ5S3D+fqUpLYhHaVwIuZgAc
GbQQxjHPT0V68TUDte3x0wHahFAEGGLAGnfgEta6ZakOMevPzJLdnFFkVmh99XSCFG+Bi9MrqxaS
s7kPgjZPAG7oAAsoPc4tIhApfDCia5MNZmHW8+s50n2K6jff7YhJtIBXlFzSnk0P2wIl1ljeWxL+
ZOaTCY7rPaZ5KC+BSEF/oehR2lrff9Rir2p/fL0Vx6YQ2BtAit9Cq0tZf8UEnyjJ4u8LUC91LOi1
mnCYE0BbVrKR/r2U3m81V4+DnMWhKgDdFPyXu4TE7OXBf7uaq+4idMeL3YVKg6vLvMj/UhNV2Jje
ezDtx3mj9aWzikLUKy6k/+pCCRxSXdz80IyAYnC0yEij00lHI1HhqUJhM+h6Zotw5fTErJBlddNb
r1e8vzb+RmAL8nh7CnrugEhHP27R7v33mvyjA3O+uFnybCNmkpMrGU+A7daKQL/JDFFVS74y2evI
3J7wBI3Z4pwSvqlnkTVfG9ZyLgpDdLwfb6gLKz2vaHWKWEAD7EYiFJBJ++8cOaDRtqTm2y7upo2y
OQTbe2e9Zt4WjYLnaOvRHCusufitOG5Lkay6E/xInWovUFGbKK8lWQ3C9/hIVbZcSsxdaMhddeqU
AIx8B9jVN9+OPStnLsIwmVrTvQggZtIvIlOZpLDOeypA58Gs6xyZICCdv6dpoMunx5CxQhBTZDOK
HwGtlbppMZZ9KSCjQfwW2GQJgSKklJjs9j1J0/x8ga3KgSbmU/Jk6XyiRW4V4QiD4ZXW+6NJeug9
eTWxy1Ft8218YKseCV3aVl6eJoPrdK9FWHjk937QLCpkGFDVzmu1E0WLDcV6psghn+UK6GPU8pJv
Fi0bbafBAjprY1NRDrFnaRH9TJ7RqLHcR1+nxQARBJvXsIXlZG0FTECKG4zC+TIji/ElyvgKOEri
2KSKCnd6384mjnJJ9MRtYBt8Zfb6bdBeeN9P0e/RbNdMyU1X6H7XN0V1FI/nJT7DXgNrdCiOHsAq
hkvCfzdRkWdq0uipPVFL4YG8T+tzLksRrY8tmhUdZGeWXxl9/AbzGdkuxAogKqTOoRbhURszvk/+
WRAwJAE4SL0cjnFMB6sqgE0/GJGhUTlrEd5/SmRM1gWUSRB486MYQe5FVIBFHqEPUkLNEDkWqn0y
+tSB+qOuv3XWY4eYuStWPz8qx/GASsULEWe77fFIkK3PzCJqs5plHyvH6dXqwFD/BFLFitRfCbdN
HnA+2z9OeABt+nHK/gEcN018TVCsw6q3pZPHdR3iWUzeoDvEgGBZwfezkK08lk22HAWNOdyamF8H
6jUvVz231vLwxvbbTcjjru9Epk+Weakr5ciMw71hODplgAktJaJkF7Irb9Ty8lJjZWkZUhGUUT0H
9NX30uS/R15iW5zdNorPxcMAi2Jw++F2dwCiB4bmvxFGIQxCUmXezidImK/HMlMXP6h7467pULtj
IbIS/jYE2BCH+8bwT8PAjDby8fYrMgJX4PCdseNGg+leRKu2+DNDnrhJSso6dsYNKO6FsfBZSKTj
tegKfAaRyy+GpqbPZoIW8XgQYFE80l2fWyLxD8IXPH6JwWKgIV9v62zH/UiW1Bp5MSkDJSIlEugN
dwVBje7iJIVq3Ddyxk8K3/rkQCp+LR8lo4/nEbXeMRjk9EsCxv0ptJ6fUwAqJ1RjKplih35iyKyE
jLxmISRmpokx68bQ3RyU7H85XLxer9FkeCLiDh/27X9r8ECFVwnfDO87lYlx6fJqx+ZEnYOmrNbT
yf+YEV+kMXncxfi7niNiqPAsZmoeH0Jey4HAXVw4rFKYNyBCE1x+OLElLycAduUVbsm3liSw5vh0
+IlSpZrzZgAXChserRviNKvo39L9UvmFlIwUMhh7yPTap4P9RImY/1PwKwGcQXY7aVv6PZHPTqs+
lzAcZRsn4Cabaqw7oQkJ/QuLwr5pxfesWq33gjPAFU/t6/YA3kmJKNOmxavo+qmzmhNRb7RPmdcP
oxmX6THs0UcwQgdPFFCQZ792AEYIHpq06O+GQMjIsN5nrmvma6AjgQGPGigfQYxz0Ux2XgitCPIM
iX/qEU5Y8+98iOn6j5gU1049fopADqafrOd/qhr1njjSDNt+Ppch21rUP3ecyG9PqqONKNQyygYg
/DuVEohWmeCC6Irq74JrYldXvCQy3XsG5CmfmWGG+EytBnU/dxqm4A0UgpUi//JrGc0nOs0dDKPF
rVnXhw1qa2u7IThR6gy8iYWztHUDhyE7T8onvmqaWONBi+NfnkJ0H+BpNXAFPh38EOGS7CbSk77V
n5la8hw+TuqxBZ6EWANW7jQje1l9VJnBYe5pgwVlokgoyNyi/dZFKwGrsfv33oqodokmWVZ4AtJW
ouGXE1CJX56UR+HJv1mQdWBnN7JOWjATCPwm3dqxkS2gh7DAAChQRgcAzcNG6KpfTI6OEPYHd6Vm
Fp7AcTVZUKRPBQopCRAjrZ3dTdEClj45Z0f5qUglfIdA6YkJOMTd7Yr0ch3r7apCrBd7f8eTYDPD
c9Fo8u2a3raAkpcrJ1kO7tqqszbOpd5J+STDctw1QlVz0reXMUsLXiFYWaYje9YiJdPQcKRUWZnX
WDECidIjGmuE/x2lbG4fVkTHIfs6kZArMRIllNXqdXx81QQ23GAWTSpmh5+nUk6ItKYWkmGBfhIG
lzk0ScagaWY91hYx834UxL0lgRTZhA0pQMnU3+OcCpsTgjCj1LUJAS5NclOnvrGOIIRfMtPER5fF
gtwwcBu4cRICrQ/tBM+ze2Jy8TzGg2eS6Ceib4DxwY9hyG88h/YQsTaBfXUPVBIFFlW1BUQAUx5r
irwhzrgonelHMWa08U1kcBCxXbHzCsDacWYEzuS2Cmsj+JETamJac/l4tpolq0G02XuXZLUSfiAF
2KZTX3Jd+3mOxsFDkItFSl6GeNGERRULnp4uvXm+Kq/W8gfyVeUzY+FGaYpdxlkCGsqmps/xuNYS
bfmeZJadMiLmXzdob7aYlhCFgiSFHrT4aV+aDu/pqniHrnbP7pgNbX6mARkuCIbE761nEBTogGDe
co0oT9t/k1oVOpUq1rOCoq9o+Yhi9tKrF2mTBo3poafo37WuUeLrP/iuhqCc1rOA5a1DVn4mrVqy
OcI9WG7Z6FwWcx9uX/4BikBiV4+bOEArKPYMOQNZnyG+NL1mlxpeVGAjNynruf9hrAq/daYYS2/f
GRsMkjX09Yqfu7gNC0bfwJ/k5/f9zuAKKsmVdJ+nP5WYEzIbvdAzuKzO6fyD7boGn7M0eI5SO9a4
cbxr1qujWnVxRJU7w8qQ79HhSrd5BxaW8CgoINVySSK7QSlRD6pk1QzyAJDqDdoKeoXYdpYXTVJm
dhRbgFyMQ+OYqENmeO5804FscQHN0omM16XFl6XWBvHI54CWIjYorkyqlszG9h/icOYnL9T3Is5L
ODm/fdPbsxHE6dA9IBtvalDU3vKngnSLqWoTi99cVrF+PFe27NItTHRTG5ymrzGaYeel7G+MOvOT
YS/Ahmnxl5TfibauOZNTYbO2y+Pk/KMPGng/pgLd+zl3Isk9c5b9EIxGuLM0Ibik0Ha9QdndkqcK
+aXcWvv5VbBOtjv0IM3wuh+TWLVxC5GbBNzaUrt3ZLf0lzoHncmJn8UplY0jFLNloHbx8BvzPkzO
v9oTSPzOwXp4wqAt8a7ls2PsJlHxkf5T/i5clgZTLpoHU3h+MKQ9yr9EC0Mkur1fXaa0abtQWPlO
diemuKHGbf6PzqAbbi/tT2SKUJ2+xbb5cO+XCgS6Ls5trMS1o6qx3QLyTI9qENj/z3tNW0k4GWIP
pCHCMc80bDHWiHHFXPTb8/zSzgkqeKjYWfTgH1HwWaZHWGURD4jFWr9zpQH1DIIFfDLuZuz0PiqZ
5LlYt/g/4Y2EfzMGrMhAHtx9MbSme6SE/y6ypsDOCGikDMbZwthJPKMkpQ310W85TSt1lT/qUzXt
y45bY1B/beP7Sflv5/HtouN7+jzOqbB5pt6gulQzisdltD3aWwiNCVgX7pBK0y/2pMZs8FnmWGRd
48rfVpuRRzCT/FX3Xqc+9JkNY6nl+Pz1QAgMTwWRFsq5t6PYggg3R6oU+h319yDymD1ARTLz0WLT
ShoW6ZU6OCO9Nj/VGW4tV06HdVa0qClNSx2w5Jdm0RVbzw8Tm+XHzlzQFWvsD1f2xBp8jFPPNdkT
53Evhk/F13Tjhdp2zRocwI6l+BQjPmpKY+i+ugXgu7udRfq2TDU1Xf5a4s+O7k6bJbXDje1EicZi
mTv1w4kUXxYt2F3yOBScivLeNCWaQo0ZqkCo0AjeWqYkkTZHHBjd7qWdOfWM6URBiRjSpTPHVH40
nPSE7NjgPIqNB77SJMogDDv2gFsn5KnDDVBrzkzR/42Byg1S7cDov6LmLAqnVxeCf/CuIYXkef+W
SOK20OOC54mUIYO2H9as5gzdhn7/Fkfpe0hQAVn+4LwOZd/PJYqi4mhh5D5vSDJd9NUvG9O4++7j
QDZDVH1TBP7nFAHsqE9rzH7fSgtRrGQQmsUKyFpuUlblutETFz5Iu2zT8IhpBIhjc9fJPOsrqqHR
bbbLFjzR04Jt8vc8qmPevvp59j5q7ayH5SXWX5ZjP7+mkhUTwAl/U/Ee8G+dzpLYDgW7PtCVKs5W
wAZxUFtSoEfcBuePrCDy0lKQWJhZc9HuyF+DRJcc4qp4wg8MWmIZXaLYTIa3sKHgVwhjjITfHQUC
mNdiblcdSDpxbqcYZUV65BSDVnfm9FCKF03NnFti/CA3zNYDyB8uIrjpW/RN6iEjAxN+t/5g1IzH
YPqSOLm0Udf1x0mb7VoVKOn9X4gWQ6x56InChAjoqg1Faeq/a5MZjwd7dAW21IerkNMcsKy0JLUF
q99+NbMdQhHL7Rj6nNXBwRnfUCRyj7ldKQl0HBJHqeJFzAonOjCEtfEcvYIcPQrYiABYNObP6k6C
NxLH73KiDdgrBkvhJrTrGZQ8Yu7mkF+7lhn4bGLvRVhWA3FKcPPAC6jjO4rMMNHEBMJtog7i5k3O
EbFM32XYPKkBnN6GPvXligdVTSBwoYyzOSxrQEI00HqIn1oSiEIHfeVVZPSCy1uS43moOpW/y4wK
hCBL0QmI9J3AS7SRlu3Hzyui89M+b0/RTVxvq9SVwukyTgEbQC8IYJdxwRBCrf8/pvxXq//Rb6AQ
9ltcR+5XDmtdW3MKCDDCHoO79jHu2aTqV24NNDjTxt58OleXzeWLU5trEh6EY9MyJDU0q8TnCWAW
tevfQ8i3JXujFnV8DShIHyXteyxBh6Q8w9RqKmUBJR7mWjz2Qev7huVUwwzlXFNcxUVzMaKd6Px4
puiVAwUIhyvloVQfzxgiA6CUZn0++T4qsyqPCESq/KrvH5az9FhcPRgu0ASbXOARHPvQi8/Xxz1q
oyYkOCGR0XeiizZfRMgph0w3fUCQC1XCaWj2h6JY1x8ZfP/Kgs3GXCRJseLJqZQkCmaaS9mGk0MG
gDal3vgqaxIF5BzfwPkCS8gK18v+i/LPWiql14Z15G5jAaBvbJ0Nea7uQzKwpd688dvJVc2o2rAN
BQYw91pJH361ZuMhfrTYj2PtNoDOBopQ+v9TicrAYhUZGleYNe3zeI0cD20bJhe/cUELMS97Q7qh
lUZaXXDQjI0ktEMBwE77I/ZISlA4ViqYaUXE4iG8TKKzwPwqcb4qJjYvRlES+PvdALS2kuET4ZIc
xdZ7m7o7c2aAvgNg2BWX8o+Hp6p+1hx2IVrc+T+zggBbRM0iKP+72L10vXK8BBCRM0pUWGzs6INW
NgDooLd6be6GrAlB46YXqaftcJ/4lAP4uDGFj9FFVpmHhw+wRbw2VON8y4OewhG5VARAhFwRJ11A
orP0S9uv1J7pQPofsIFjaNQNLDOt2yRvQGXQSPu/9TOgnGp4hU79Pex2PhkIhGeVtHQ19CIoJU/n
qlAGDMG+J/EIDxrls+x3tRyBsiMlYdFeiwdaR3u15sva1Q3B7uHwUHmu2IYuP4fe4Lqy9/QXkeFT
c5mzkZV4/CBX763jbOgikgp+pcmKM62kzKRwRmnfx6cBsbZSyPksR9xN9BJ7JpGceo77/FkNJuoZ
8X5ugJTfh12eASF5QGyCfPckoBDX2Y9yNp1pq314mKZQfrzGIiDGEjDCtY37m8X/AmoV0xAGScBC
EkrF3LhCAZ9LZ/TvNmeY8hbWjsc3c0xcK0+6dmnEyLNq9PVxJu6bHDg/1sdX2Ql7izeeOO/5IuxW
61+CxncVE+Ph0/hFpwoJ3fp7Qeuzgna0jX2ufszd4L57ajyL9LzGylDyHfTWGwsHXVmqLqWlYSz6
xs8mHwCnc4ku27YpF5mqTxnRyEefPCkBYlYuJocAgorX8D5yn3Nq4RE/KvCSR9mDgZ2dg8LocEz1
RsAuCj2q4YuHLFPoEFJEzGBSKxziDsvrYUrMhTigIx9ehPNjW/dI6QDhD/ZbCHWUFjohq1q+15Y5
tM4qSR2cwqZy10XA37CKiUFmLjnthl1wag4qI5jvyU6MOapf5UjZGfFNlIkLkahifzAK4C1TjTZy
AjvDHz4Jt7KejD97ABSPxxaEBCVPPPRXHI54cjm8/RhfJNlxqt0PRlECHdBFDTiv1I1T9+992G/4
GWdOK2E8l4GFn25USi+xXZv5aF8cctOqND9y97MaUgm9dZdaTQksR5K9yqrxf99X8hVxp9VLi3xO
sJATWp0IGziRSEYcD/xdfbjhuavq9p/nfN9zP3YSpyIT4yjPLPdOyoGDFIMQ0mveF4PR+FLWlVn0
JKLgNM/FfCupxWWiruxsfSkUJeJlGJ0BSTEIwviy7tvcVtgaT4ccSTPBHW8n/ADg1hgXzOi15qAR
QDBHtXXCJA68PPBiIgAGPhwfFyoIo0aiJG7STuPWtvOE+1M2AqbucgtzYmL6ApSNWq82uK0Jh7Hm
8KDrG3Zx+e9X4TGueyROKrue+6bsR+71plHLN4ZnDQdn1YkPj/tHir25xiKO28mlRTl8/PVt0rMh
cEPMPgaRqwGrCPHX8Ju7R62xzJc33SPBwIFcGll+lBHVCkRMxKPcohsxnuYe6I1D2nHWbbvxT0l5
BDIvB2wu/XvmvfMkeK/D1qxflRhWYZmeC3klBOLngga9xCzKORJZoCrYFTlzWSyPRjT1avlkDzg6
S8jMAfxDZwnCapvJaqClofXGfYQv3wRF2lJCSYXCSY6ZOPEtZ7vh0E+SA6ruBQLDU0HCKjK+zSav
Asg69KNywGNRbREgW7aL1G1eUIErl8FO7O+EAJ2Not25AmOxy8+tWTy4RIiTb8/e+2r5LMD/kVau
fcZM8AJGFW8va8ePad1KQuUR77c+scwagn76S9/oIAUZwg3rmWSWDiqrn1wTF7m+16Q+DFTYA1KW
ls2X2GqweFOVlGlOQAWCp03e4emcfZj97k4rxxGXElFtBIsKGO2FcyIr9RqbHZBjP1PdWSswRi6Y
XbHniXLYiqDORPOw7Y4c49Ge8E93V2+aAGCQ6AIcK0PLS18wIFBEZdVyk/I9kIFhRcQzrncHoJAi
CicsqNyE5BZ+f6FkaVl+j2qNbf3T5kOBrh7mC8OyKb2ylxtJGjJZglfs3by+f0V9YQyxu/+rBayC
dfXKCOEh1lSzN1p4yoPyy5mkAnVZ3D3Jnj2rvu3jHzKYyUbRdT/e8uovCjs1CRsOdebebDss+aTe
gfFq/uQqOl8XwmxNjJq4JWFDlzY5P+9b/ojVKnhWGXmfS1HWHo0DZKwY6i8wxOWEAl+elqM0WCCI
6KJiW2vARxzvMDm5ZY1tT4SIKJzy/ECA75FTbNkUPWRYwXlGw4lQ0g1G/jnUURxpvSVWcpaWLsah
eyjbe/KM4fF0IObulvUSJijS+B/AI7QeeZuqo07iLccv+/COa9cS2mFPaIvw/E49yq13yHiQA7zc
AwSk8WfHn/OAZbhGyZ0EUWintmfMDQi3FY0o13iN06hvRjhyXgP16VReAS1qCTI0cLtdGjOyaKmv
tPspjgK+x58+6k5kPBIaRwmYA6Z+vXu4kXZeevx46v+wr/OXVFl4Bn3xYkV7Ye/sMt44+2XhFfdj
AO0GA5x7t2vl5Prs+eXOi9cgS9a4vjyG2wSM7qZLklZUtYKXXRzMqrjmuwLkC+YBL33bfhohP0IR
GuR38TgsENg97qrzPPj2p4KsZmQFNBoDax4qDWVXZG8heR/mQz8dKV0+LsTaXl4ZfzX/hMGFVEhw
ZIaxXNzthDV4AZWVpHtv1jl4VITOvrClmGqMVr05aS/hbqeA9b2MV9egniXeD8bY9fwbgUqnIzvk
ZvC3uVett0m2vucrdh24mfRT0F2bCZwiCegLL5BOdrUe+HheUexVmBJEQ6DJj5IXVRN+vOTt3fua
USOy5w6x7i/oyi0AgYOOJqmFGLCdNFeH3dq6l0ZbiiYTQDJzIrigFgvnZgN8qLL2GyovURCGFVBr
LUmHwl074QrFkf4m/xUXziqLxsJ51/pvOVmEQoxBAJ8IYZ2Jw+QtYka82AtCdIaUwRahaRMjaOsa
RBWcd2MOFkUAGVMgaV3WBqx02lyxwrKAmFyAdFQrpfu7lLOG/TMxBYTIHUvRT4jFyfFf2l05Rxy1
TQn/YXy0E9zDaO1NUAEYW0saF/A1ijxerGyNraG+sbe/ZBt/PDiMBdopncbmRoWmeI+xpFOj3mw+
x8u1Qg04cDQAqWCLGqRXiGvP62nIzkjnf4SXbnsPGYeHBRfz6uD9uR++9LFp6k6ru+aVMoGcZh1D
9DjoqSlChqt2mbHPwd7lN033lEz/fbIXQimlMYHY2jzaBvskIleTrYt3J3q8eYS2Vx1ftTuFZCGb
eFpGg5l2bYFBl8Mxmr/8HQCSZ5gecyKcrnPpZ9jCtJD0++W24dzeBpMTPtwpD7p4ueT30gWQzKR6
cwwvFbqXA/taG96ja1ipXUSHBrQ31G5U5GTGpjyBlY4eW+kTH37eyMeNDj09fENjEzJRySiefej0
aTMuFUQ8xSCseDcpfFftGOwXYYinhiovC0e63UxbO4n9Zv0S5/NYu26dyXLXKzdx3yqf9UhYXiJd
OWrRPN4M3zF7jiaF92q8LvSf4I9N0d4D+V/O4GTAEaqivHJU6tDB7N9ltUrRcITwIvvbGvG7iWYI
fWtHVflp0EaxJWqNaEqsgGEqRnOY1ZiRVOmBSkesbGCtVTO0FyQyQN0zhgrNiM1XafSmVMByGi2O
2omYeG2JTlm7OMkiOQTZEYR6Ksj+YQ8huQOKxk0hqvXGWuXarUGSw5DoNRHo8mnh3dVNwseFEQ55
KPvr8uOwv/az2FRR1khLwt8lDxtog6S0gxPkKbAs3Mc/MJkBxg9Ymun/IiwmU63IQSBtDW3Tn5bN
NBq/w7knyaHBGpsCoegIYorZWilR1AWKjLPJ1CFbF+H6nygSwx7vrdqfTFfrnARl2QJD28/Xs4Qr
q8Kjyu+CYJRjrBnz/pnRqpS+dlbWK2oQpHKZB2O6vfrYYX4JOFka9SghWc4lN4s8fJvR/Pitr0Jq
0lCAHGJn1few7xM2kSe5zM7Z2V/Ricf1AMJke7jT7ZRmlFw86QPLKZ5KOX8lcsS5cjf2A6gO+E1B
9CVIvHxiwl8mOPlJ3wIFyVxVLctt3d8yJzd0G3okxUoMwapPS0wTOjzLzpfRyoSp4KV3PbKVaMqm
ozDEiV1698kQQ0LUUmFeJVZHdTzcnGGDOrek8tAQEfPmRaUwWkCzY+iM/5giU+MnjemyqkURpsB7
hbVTuFabWnA41jfJrik8g4kPz977tcZsnz5WBY6s6HvAEqaeaPHBNx9ktiKaNBPL2yau2Ymsf4+k
g3hY1MG6OcvAL9kJiGLn31oFhUI+gnhi7dFKfURqIPTZ441e2IirqpEkQ6C/Yw9himqQvN6XcQbk
+SCAMSa4p/oa9PtwdU2avcIzgF1XJ8RIlztsRDjkAsGo36NszV1/zblyCEQ4NnlJNQKI7DRnSOLH
v8Lk/iRMxnx71uS7TlAGaXh7kJfvp0/94f6bUbo/6lwHOEUCGbOjpi0uTKdribzRe7tyx0jxsUY7
x3ia8+Q9Qj8ZAwSJ5KwKqUwuR46jQuV0gLbbppVI+mMRp6TJZ1KbkLPgyP3CbSRyGNCBbD4D7cUh
GECzFFRlxAhR/ieGwEI+dIqkrjQasKtIQv448vTMQCQH7OsqGZcfDkPehkW5ldN8GHOekvHpreuR
OgofKjPlz50Srtc+fPy9qi8XYanei8b6vQQlsvDP5FnRMg5nsp4CEMSN/N4hBFXswu+hlZe8nM0b
KGvhY85tV2gV8akaUzNkCle0VsqfUbB6pCQWyC+AAO5sdvxiuihgf2Afa6LXaic3AXiJc1b/EIHR
FI57j7W5Yo+f9fEwrNrkSFzbkvLCz4sosd6t9JgJSm2uSlg5OLhRnQVqtXlyFAFOAT4Gho7yob+e
5a3tVbBTLzMf2GM1oohXUynbfADG0wxgKLcqvUwb45N4wLp/DQyVc0ZqaP6XT6vSXITY2OSdRMCq
Ld2MzOfEqjdAufGQbmYVPfdL9p7t2JfwTWz1nQH+Co7bg0M+Fr57X+tXHHPHYy74vzhkFFMCpR1+
krBo4sx3vv05pRXnaERJfp/Ooy7PTmc6OVb9llJAW5r/dYebJEsCpQimERG7mAcjutk27NATOs3o
Kpx4/RjSDSJV9wwlAOv/yLk29nl3DR0xo17FTFTR3GjZM7bANZR36Jzd1QOfIaVSoHXq4V6bU2zo
mtJtzuD1IzeI5gdMbjY7u5gg3DF+QR1FY/YSU+tARfnbcEX88iakV9zi/wNAvxVHTT9I9jL7g5eF
7P4OagfHnlx0ATZ5Gob8dWUKVAxH7BC+CWpRxRWnK4LEunZxZJ38hSTt1OPGmRT8YaUQ+r1xrSkA
F3bNuJp+EGzKJY+f21CDCVNIGZ6l5F+uERE0lJSIeNjgh7dYzbxZnyBZQnytITMBbYkW87ZuaGAv
IxasPNvfjEbtYKhB5Jn1UmgbhBXmqTTcG4HlbbNFjGYVbTZ/ywZ5iI6f1Jay48MHMI1alQO8dS34
NZvWKOnM/Gfdo5mdbWYamt4xAgo/Ohk4vNUJ0CHzaxqR8/eaW7UWUDIGh8RxHFJhw8qvZcCcN9kV
Cj4L5sBQ8UUKC/RTGWXV91RAOAz7H26VfgSeiQ8PZnKa9SQZhcS9V+B5rwvWemERfD1wzeGmbAWr
RzKqaRUveDu1Zq51+pltNDA68xYLEOtV09mimALL/nPshwb6Txj4+a5zRRbJeMOeT1gzoEXsCOsf
F5wMnHYyAD6/twhM6Axh/FxFw01VadgjxTzepNPDTTmOi5lC/rH5c7vVwnvlPv6UC0hA7OqFYrdo
uv58TSYNIBUO9SLL81wrlQzHdMqf0iKiUW8WKulcWx63gWaV0lDPbC55RyToEwy5EUiG+rhWs3ae
lpgInWOgTDdhsgnOJ4tA5GYjnu+MJBsMHp4II1GA1dcs8UruhA5hQVribomaWC1bxH0epTsVNC96
jbn9vO2HLecKXQz4UX+8TEcA0MlN17WHSrlXguXiXBx42uwo804N9wfWIwoZ9koSWEkj1KsrVLDH
d81+p/9hvdDkhDzlQhaKG+KUIMqFlcGpKUJJpq+NowS74B8GysOgOl9dAEG2emJLELcC8RtLCs+o
BeMV8+oXD5RLlvbCpDhSMldSiaWxLpBFZkW/HDL2FKvLT/G5Xs1hEoamDWF1Q6tFQfH0DsEEcjSt
sdNwzBlugicnjTUUAcrKZ6ZAIaFL3bsYeFwQOTbKn0L90GRsp4vqkZD+Lr8MsHcNZWnWVNMDIIB7
pg4FxmkqxydNn4p1I0nyYCFMLUckINUIYNfCuKT+suhQ2sABalzcv3rNy5TEH06eerJskGRscwWy
hlPSQA3tR2NmcFG/kTEqb2ABqFM7/plYw0CNvhorgaSW0vCP0EtWPKHOBtk3A8kujveBVOZavMSS
JINZlLS/Bej9hi1vHneBcIMh6pd0zG3ZbOwzuYMEbgU7IOmsIYXLdHSZG7xU2MroPX4eIisegMQy
jRz4JbteZVWZGDI389avY+AvAwm5+1gojej7bZ+aNe+5uZdHNpxX3dTL8Fl/yRpUWEkyxNC+Hyws
OISpdf7uuzirhKt4vDJ1gJ3IChD/e1DiAbrQkYGw+DbchD34+qs9rdsiNlJDG89CwSOBtHzX6BYd
AiWdve25WROGbGyHNEijlsd8V8UkoecSXQU+PVaGHbtVfbVXXWb4wg+JqOqdZIxBzeOVnVa3aXkT
FiHLDF8d2VCJ8TR88yfOf7NrEXpUlJkiFQrv3t9wWOXxuNcXEZDCATCy3I+7qi9SOayGoK7Jmv0p
uomIR9DZZS3L3i0OZBOeaAd9bn5L/UMmpkVpP1o0S+Kp5l7sFcbP78d+0JXLdpfQfvE6iwpodsnA
uXPrT4vfO0ucInFGF0fs8q8US9H0kaaOOa8iV2RD/xBIJxBy13nsEYeTodK8UA9wE8sao9kj7/XI
FzrW7y9c5GsWGA/XYrXH3/AQQwIpHJa8Y7EGXomeLAX6Z3a1ypM336Mt1397KE7c5R+MG717/XbY
Kwf3EOAtPPuPqY3JbJRKg1UD1wXV9X6kmoThcA02QsiEsQKlg20P5uYo6kUoY3y/fT1oXZe/DYNt
g+iJDnxya8+14e3HqoWOb5JnDili2y/5jXt1UbC2p5B9y5T8v3G+vUVL6mfyCmm8NxPC6wM6j0IB
fbFTkIMQCxaF06tivGdQV4AZ3oISMo9ANddNPaG+Jb1d17YrFv0cBUpUN1UgWbcEoAMZlpfBJ4m1
UyCAGmZwAWKtp+oDgtC0TANrGM6rUdJ9ZfXT/Z0cGiKYN0IpPIh3H5RdptTphrNmdG654YaOI6IG
lliOfdJG7SPuowoc/A+AgbJxlSDZtT3iEaN7icYqLDnyZCSBIl1mOIv2wnGUWG1oPdTCoCleHsyZ
+Ny+awYlgBXjtjTWg3Oacwus3RNtmdb46VK9jlo0xnN1jHZKnLsG2MvMOL+U+Z0LhX2Aw68sosKg
fn4Jtu8+hrmufMLUjwpi+9oVHokFsIlQxDPKNmbxrHZPyErw9Gvd7ukjYz62EDDkXMII3JO0eN8Z
sYWg3q1We7UCwof0tg8rhpJYqNPFQRA8cO6yWd2YlgZ1U65o4amEDtofXRFfdfdNhT54HHIPjSOD
JGB+DsS62eu0zQhiksWXE/HGn8utlXk2tnP2J3SqTzFRZW8yqdIW2zWW7mGnMXs/Jal8mcRHp8p9
31df+zyvev8sMhcXFuPgCCNrJJ5EKjSW9eGuj7IwIxQ+zRuA5KlOHL1FqSCUDySEn1b73w34oX2M
9J40+e2AShXPd15YaP8c3ExpB0mnGXAkZ5dJZMwyw8f69mAjKX7xBa2DvShyQ7fKO8NyhBuUTzea
xeFub/L1C5edj+6r6bKrOLp9IrAxNIAywWlGdc1UWXsKxzh8EjugUfyO5WkSeQnvlPKU9h1Svwgm
2wWwf0Wom5U7irHBs7B/vPr2ccytm359mhOgoYUcT1gH0L2H0yGLiqoyn2i4wIgcI5mCTOVpRM7z
TsDa5gM5KvaTCvqL5wftCxAMcMr3qX2+lD1IIhuX26a8shU/eseoTBoetxIfzipsVLqV+mLunqk4
NRiuaDQhhM8CG8+JWAn86hkyDAEZcbVSDHHbeRcXhMSoAl23KQL+p9fdjwqlUoQNgWCFRS4BrAsv
EBOoD61Vz+R8YVF/HgCfIwwwIeeEa2PHh9nqV/QzQZ8hFeheac4J2gYZEy01QeC2KtZw9i06x4D7
PFgr8mYACOMlZ2l/tsntyoPLk99ZGur/fHls0nRvIEUi9+P/cfWVdcjfIcsqTVDf/REuRuW7HviZ
or8vYbIzDTjZeaDzkfJvrE738+27iHK4kDCsOMFo/PC+ocu78e58iV89Cc1kZIWk7bGTmLb4Izys
db9lPRNJrKw4SZ33WkEIakDQR6AoMLxp/qj+vkY0fojBXVzFPDCNQX5JPmgNGr344oAy5BDHS0cs
W4wGVxjnQl0bIZXTd0XAOprJYYn9ecYFXKVrMakTzamu8u/rDkk1S9y/RSdtW+7k5EoiFDk6t9ev
9c7YoO0THOwPP/MEahyS1xG6+oApd/SFzwsuRqJWnDzIFuf5JaP4/RZI4AwuBGGQfy2TXbm2WI6t
eAujPGKqQDk70RZu5/6HzyOWDgzDN2WMOlXHTXe7CrCv3y8IxUk/xiTrY2NjmtXj7tzb7+UaEd3/
2bOR9dkvvw++nylt4jg3SFglApLRkvSEu9tfl8bL7nCHxz5lCDgZMPC2Y4q9jrlU88+RZ4NEmG26
CGek9T7cB0LtS/+F3u7Nxivsa+HAXjq41lg0IrDBVxhRPnfbN9DiTdWXloSqdc+6Qzeo8c1MOBlg
pRFBDTYGn4c+ryMLBSM/9f181QqVjezp/IEtStDPOfmFdE50eIcRsDaDLZiFx/ZjnLv9/aS50Ypi
CzTZs/bsX8ZTiQCmg+xayyx9+Afw606DDLVezG3gq4JE4QT3U3g0YwDitOZIXDyUliL2JheB/CJP
j4taoxdNBbpJlqd5H7YKpDh1CnC1uO8x11kliqu7/2wO+M3BekOH6X1zCfWGqbGEKtsEsPyPZPyc
LhP2wVD6+g78ewx58GtchfMFukHd8D9o2xLGYrNA7GQWpwJ+Lq6SpIja7PN3XByGsMxRR/0CthdB
YlfHh3wv9OiNkH5FaQXEYo/VeCoSHVhC8Qd5XFMyneEvXZ/N/SJxIcFU4Zl3PsP1cquUSwbjsCPX
unrrKSBfuZ4cl0r0wjwCfeOYXjsuyVtAOw6lRuIRXzofp7anoz1sf0W7+DaLVofqOMljs3tzzDVe
mf+Zb43+WPMi3s8xZQPl41OByrQgQRcfX/5pDZWxtGeH8lwKzeTEVXytqhRN+PCwIs83Cqslbbry
d27gMts1kozBfieog8HC8thYxZYQu4L3IlMHhTFs0Lf4R76kaEMY78pGnOnwgSpX4LeGoyzwxa0+
89zP9luIrkbLvu0RFV5F1ezHGuycnOmGMHupO/MOF+Vc/gEoE1uwtekAp4un3pbZ38MVG426l6vI
9803CvI1XbazrKuuNPRgWDCl+xzlMPN81ix4lCTlbgDSiuIxv8BCmVFSP/AnjryjHS190EtZZdIn
qL0kd6yO9wp6y2eKzvyOB+0sBRH/dYr5+IGejomBbiK+C+w7MV40pTwnZWzItC98CLrzs6VcJ2cg
j6GjHI6vctEg++U0vdaOrqdjS8mlXBZ2E/4fPTZPUdV5J0gJJ4ZyQUg8TgQpx4iPYiDNoT5+qtPE
txj4373lkdHjtks0CH7VUhYsccHyXZpqTW7VuuPdrnWA6ag8Aub4vNuv+GjzlweQqLEbt6sUUHrR
YoEjCqXNC3VtkrVdz5+8goYAmi5AEK0py9v4kVyoBk131Gp5Q2VyF5iNtGrfcl4bmROu9LSX+XWl
j1xYDA+dwhWNgtRQc6Xa4+HLph6q1lM59O3uGtDScQlSmlcM0YXkS3wPohGxj3g8vHHb2pPjA5bs
YUH5ACc/gSbV3eHH4QoVzZphXJbDPlMEZhxX4hCCz19XObmv7EKt73ZJ/6JwPzVRH9Fo+HBJIg/w
6IlsO2GEtSwLICpyXXOfo22gdo4IXPksfKfFb+ctNXZ2g4ZzmRzQ9FMn3oMkpqaBRlGYZ/7qyQfV
C3E7H244QZbhI1jF8FMja6u5QOYV4E9CKhSX37jlHHEw8mmnb3wd1OBV9hVG8K8bfF6/mtvjb3Mu
tcRk3nd0ktwMW6hOMDWWJTPMsI5NV2CmI52mXX1yJRL98t6kRPxXuLpMxUFYH8LIujhdAib9WsQI
dL1p+AMhxz6ZB2tLR2pQ22C92gJ9PZFPNavuSE1GfQ/bW9eXpGtExszxVMkkaOnXpKbQfUIzM3ie
TDh0L5NX7MpIJY5e1f3JB4rvdaxphVSJAiwRnfMeYdz+A4OFtblpYuQAFlS3bbU8dCsJfS2E93pc
5O7I8GiwyFm5nxF976coXmNlcSml+T8M+Pr41NzBFnRoianLzyHlXh+NcTnxe1BxgqxeazFzOVQP
qfE3RTThHvCq1fY1RlQOiVHUvWXSbTS1wbAFdhyIWwBZFijDDPHh0V9oIHVc6W9LVWUa/PTE74z+
3o1fEiFpJ39vOCTaMc/XkkJ1O4PybbES5hkx1XNQSo6ygbdnetobPs1I5kfyM1a4ccGNHznM9ssp
eCCmLcSN9XV2SWMji3pUzQkrc+yZ6SQhalr1smPAarNx9/m0saALQWYX8x44Ur42pPX9ycwH+ijw
vyTLXowqxo5eU86k06+kjG8yA/5ucNPhpKOzXKyjJBr+DVB8zO+L1UFFaasX8b/eqNx3aMCgoggN
/Te4KYJTCB1zxVHFa38aznpRZCYV6HwzlaTTNmJPwKix1KsV3GPDnHniQiBnNdgYKtzxIoXv1NqF
Uid3BV8ix5W5MpKYrmzS81BkNj0kmgsLRv5T6nZ1E+d05L7MbZpZi42OifnppzuvLlMwxWHs0Iu1
LC5TKNt5sH6uXnfXElu4tiJnNBLlQlFkMvjJNhz21YTsRBMaNlDCu58LfaCRI0Q/0wGknQ9/ldj+
GuS3qQcfa3RMCkMjiAPA4NvqXFVAoOS1H/DRKrXH5F/2Yy1PgEig+q0DKcKbW4a0zwZOreTkdtqq
i6yoPBivUyeS2wLyk9kZe9R0ejCJAqw7s08MJRRb+V1vABdQE238pIc3g0H6kw4/OVMPUljomPUY
30TVDhCB1tRIG/Urt0YJM3rl7hmojmq5tse4scpDuNg9RafsA0/VYDfivTiASy9dXKqhSMHxA0WA
abZAy3PfyOQNZXozLihUSlHY8FJzdfZUhnskLbjDMe3RyyXQHzaCyEO2WHM5tUSoT4BlzDI6WP+F
Hyb+S+t7rwQbcuMCPNrrYW4lYcgq+u9sRF1JepWhyh6uGI9GuQ1xE+ydtZxWVU84xcJ3ZtJDTbo3
hQTOFC2UJ0g1txEK6gIU1Figkq5Jp5mncM/knwjMhpTaFkfxxn21scakD5NMGYTxrPt+peoowX18
Kzw/8X/Br4Pv/rNiIDckfGSX07LP7i9+POlNqI7cXmd9/S4s1z9tJUrBiB7dMtG32Mc244mHeVoa
9CxEcL99rG/mdZuZVhFayOJ51DC6aSkndQIaV1FAL2PJ7C4l6nO4Qpnp5keMR8ZzkQhOYNHD4bGM
9gcZ92GlbB22KMVOSelnvJX6YoScoErjJPmD5xnWjFc7rJ7jcLxQdvpVfTgtVH4GVc3h1FUqbuTE
slKNuUdLLdS0sfAbsx89ug5mVV2a1ucXqylWR5ZPtlzi1LXfS54wfGKByCXOwjVUebaNlUy9WxAL
QmIpjaLwsdKYir0Y5/sU3o/YU3vM4+pMd5C9/cJSmPI9Tt0qvVSV9EvIYG0YmFnFg32NyNcHZYt3
UdUBoJWLuxbk/jP42Iq5QzSDq4QjNND7YuvxSTtUTesxeYI39wv6+63adNMIA62UJWlYXYa3x437
N0vHwGNLPC7jNA8DxA5VE7EMKcLKW/IcGz+kuKv89I3Y9BAcP7ZVCWUuf+tZgRJvagqG3u/SS4cp
ybjvZ41/6Yyqmr43Mmu0BE12sZehnYvEFTOX5jzu7ZrPFcSrlOTKBjuLoqNlcOA/HYbipEF7bpVx
8lRTiwT4VQP0zYaifdqsPnJ9AnIfoThnxVnngeIQC+trGcsmQgPi1JAH0OVlcsOuW2ZAJfoiCj7y
oiES4YxjMzy5PHOfcX4kEbE6SW5xbefo9ytTTZKLyZk/D2t1wQD75FYGJXCN3lm1mewfTaprZyXl
EsQyLYQfFH59XpVOHODq0Sb8TipFqSj3zwsY+HXoOvhpka7d47riWUOGyLJyFfAs70EBnSKiruJf
+I6PPr6mpkUWMClrxgr1jTZVaSC9zrAyG0y9CSpdjZFJP4CoPh4TuvqtHNvU6/WATBv8feBKvtqh
cuantaqpT8uxORHf4CFvqwmm6ABs9mNsiHrpF/aKhqBwZwxt+5mkptDxvHlBChxDX16TFKc2eZZ0
43z0Ief22MgUHnjbc7c6JIupHPP6nI/jUbTql4m3uRMInbiXDaqbZOMfrKefbqSE0XM16Gtm+PYy
VJ1yW5U2wFEVZUh+YcbBwA/1O0X1oWyypfd1vlobOv/8fX8UOQtZP7m4hpvHvRJjcUJFMS4XTe7n
g6Ets/qfgazLT4nXNcxpn3U7GjpLL4NWj/YQ9TsuOEioGTqyvZIkarK92Q+EbnlpuLCY5icPMvin
u4maWIDUzuoPD6UzkohosdIJFaUUNMOOqKh6DQRwMBlt5D44G4wlIbkLgM0m4qjX1AhCebB5QDII
Iio5wTQ6B7dq8n0TlAa00/g+Z+haWENwTVYDC4CdqISwTkPHKBeUf3O8xRQGDUWj8XFjNqGoGrSY
2rKrlazrEGlJRrZhzvHrXmheUTTreyALXgK4PgY7Lg03cMuPkJSxuGF12X9AZJeRvgzg+1rvFHDO
Z12xsukTRKwgeTGt81UUbbODgrCaoTj/j1yDT9DMWoxNuYnIVXnyZZw9gFw3kRdg2b7YxVWIOBGt
IjJUq7iInbWX1zBKA7NaK8aa7XUMqiYIWlGr+661xR060n6UMO1StJfJCxHKXMhV9dS4GgWq4Szs
hJHVQa3J9RLktRYjIMpnfJx2b5wl2Hf076MzzgA4fm/XAr2s4YMaz1vlfZaOsQYsO3ygJslKEuj7
SDIKAf04nWOkhsf/k7JqLinJqEniKRDlwLUMrsKEACE6ypc8bsM445H0/LDMKSCqW4XPtmMpk7XF
DkzgVb7uacQ4/6GRD1BoKZzCmNMSTdmyoKLDsgQd1jwcjFwys3mFNFEf1PTJhzDq8BBrgGEbBDjg
S+oKq1G/CUry/SjSkimBPIYK3BMo/RuWVbWn2ud+x1P6C1WBRXT0/UYK6zhStM4f6DqyhbMgNqbN
ZMQLVs2ICaLArx+2Ju/mjK/Va9Q/K+FcB3MBrbVfW67C9Pd0ItyoKV/Aw5OFvdk5hhmyvCcIVu8f
Eq28DaWr4tHaQ2egRtl0PyzPu21v1BFG000GCKyUMNCuUimwyz3+ENwyWrhYmjYZr+LwKYkBqz/D
6vfVeIeq60p8Wy4FI8PrRWhuJpsV6fDSQn7iC62294HX0xOhmppponMquTQsGhWmgPChod7CvAWy
9QLD1qkaO8HGxkZDHmqq4ACB4ZaHI3WE9wv23Qb2lW2pZu7te0Ge8Pc7ydcSmjgQvaWii+/NQMn/
IP9LFvujzRr/uDfIGNvd1t1pN1p6eOc16JDOtSSz2IU70277JTKXIqiGS90WGBiEh5tdwjBUnhw+
G9XNlF0/6dZgCPrOSqO6SLdXtDnc1X8dHJAT1MAVkvxahzJ0aw3xuzTGfyMtG7F0RpWjNMq7htPP
QoTMXKadZJTJJYJK1oTIeXjd2Mexvf9m5NIZGT+EjbomcKqR3WYKBuWHX/vsD0eyg97tnCtnqmWA
7/GwEjMj2i1tDLKBCL0aRm2WC3zc62SJbwdJdXe4Li2jRpfYNd2EzM5n2M6CDtd9Th3wnYBwNAxd
K/j4WnJb+2p2JO6LM1YeRPq5829PITPrW7hbVN2WDm/uahoONCKNIvOSDMCx0B9eNZCTVNxGSyQz
r1tqJEAivaIoazjaEaGNlV6s+5zGPO+3VN/DYVlyBrcD9zlhnlpV7xWeQuD9bRsOmzLCTnag5ai3
dzNXkcvkykehEIwl/IWAZoDvLNOKAeSssdlei8r0QZHQsmB+UN5QUYCX1MdHawPZFcwUZHQWhfT0
F9R0YRvaYozLeOv+4DO5bcIIMXolUpXjjBIN76E5wVtuMGTEk9HTT+eYrfcZc8g2iJ4pd5al67Pc
Bf8IdZmoBRyuH/6xFzLOd6AYyk+6DBkpzDqfPLRXZw+tKtBDO9CBdj08sMy58ISME3uOJJEjYpM+
o6K9hb+PMf/L7jdQcOTV8/lXEoWQfhzDSsOiLMPMutIZYGr4Kk4PuonaOGKQqX+pNhC2SSChuz/d
k+tIjcwIZRFkq9pBM0X2sK+L2brNgCWOlyVvsjFgKNAlxXrnqFNZmQElnsJNFXiE4K+Y6MAsOIH4
IOnqEfQKpaM3xc0zfigZ9kUnCkOhPkKAuwMRrqRvOhXiYxPtiE3C7fEeddl2udwo9qkAw+Df0R7V
gwFeOSNs3qx3Z/VF9seLwHf5b0lGWWF0oJ6djpMWhTQlauva5n96LcGXyJFyu4F2wPwNOiBgsKAs
2wK9zo2N9mdmWnpaMTYl9RBTEwn+VcdeG31DjfdNsBwEmqp6fm6nT6NXDTFlX3a44FmZV4nMuuGJ
3zBoYOqUIZurVZmBTJo1UqxLXgb0LQFO/0fXcG2mjLFqKoa3gkpPrixXk0u7QsGDc1POhotbFIOs
FdLHI5L0BLBM3oFOJ/ZBGi30rj7vniojmLNQLsgrBYo6nIFRmWG6F3pbhR76lZ25z1gMHbEPLYtT
bShYvt3hjpcgu/MLmAEGv4MicKa/K+UWsQjg/Cg5jlxXobs4/qSbaSuvegBWYP53ikOtNHqh1+UU
cVeqj/f3FQf9gdF7UQSGREY3UxkdQwtZp1x7fX1VAwcgCjs9TXE8BoVUMW6grRmA1uHCSJ4rhil6
TK1mi0eFr5JtZbfNWSR3k4s1MjvZLqTM4ZayvMzFXoiyJQU73GSEDnVtayJ/FwciwQc0Dog/zVB2
yTtaAMV3Qpq1ZEY3Adcsa8+Vx2Xw3hpwR5hpWhEuTglGJGeThDRL2CKxstl5ajGp6JmouTKoxE0R
cAjdANhd/rHN3S1794zptMN5hyWuTsJf/y98kH1jGLoSLo/wyFpM4VZbRnEBWrYWeoYOtdpcvbxr
7tynawkvFYoOsGlHLYbCE6Npi1GzwQSEDPvEeh5HtLsU3EX0ny/yMTOQeAqa8gDhf0HznYT+bU4h
Q1DfMtv1RX9/Od28d751XO2DXt8RDKMQPUMEMtgb39i2d+FVU6KTXImyTj+Tx3FdurA0E2jqmQ9s
EWJer7VBRri2CPbpkt5Kwm+EgxaNmlXJ5YBJgN6HUCGi7JpA1Rrzwa0geSx/Q5l2FAiMmhlFFseD
bFVxWZIKVxQMUIvR6UBAu8LCub1tbJ8JrzhfkZTFaRYEu4TdsyaUmt/bcV27UaHscrWGGs2ViVwX
vp9HspqCpCXvSPl81Ecoz5VbfV59166+B9Q6+MKB6HXsgqqiAlHH9m5aAgzAgwgLABHmXw0rptD8
IvztnDBEdTWWKK4zYj4l1bVZ1FGEGJdnjxR4qGZHf+i8o49heJiHwIVS8CDteQwTAjvFoyZkO28D
D7A/3WiW6SisXEV2/ZGE2cWaVYHhUjwnIZ4r/py0LBQGZHsShOYqEdisaFiJuLgDJhdepRsb+z/4
Dxg1N+fDW+wQj5ZiBs/tn7ufeJi+9ItsW7QdAac1/A0eo9yv+Nq1IZMKP4j7p876C/vZgDXgQzj8
xNOYnuMPUztDxWmkbJu+Rm3fbRly8rM7eYqA8ZDFh2rCBEOfNn1kBb4GEx0ZLFRYIgyP1FefHSbu
sh0a3e2KqZo7i0ZbY10W19kYJfnZARG3c9YoiHzBtGZ6G0Edx1wdkzphUPV7bpxht9GDV3poZMs6
nFbWwrpR1Gh6NldlPRRVZF4wZ9jkYw69dzkBAhNi6xc8vhPKZIW4qhadXbuRo97y+5t1gmFZ0rir
D2w8R2K2i1BdFWzKcBssVX5/Rqn6knpV7lKV339Io7hiKIz+o4UnFOhHew59NRX3/CR7v1WlMa0N
w6Px0ztIKijppd/4++XfvjHJSwtLxsLwHGZZeQClW/GjEpW++/putltPNCGAW1fkGloBXUVQMvQC
dcfMaj2hCCPnwptGh+ZQ51mEuoIVc7qOCDr4MU5yfJuxHUxZsEMM0yuIDFum3ZnARijE1JuFGcVu
zqou5ER++mwMI3nNRDM285lJYf7XHq1jMSZvDMNx2rw5a13rzvgCvQQ7LxwRytDSwNkScAHAmsVF
b1xUVRv3apHO9qVaLPgER8XT8hDXA4f/VsPq8uW5SAoLgn5S3bGuY2MuqEsK7YbrOTXJ5Z8hw9Mf
S5bi5o1tmaKi79/sn9/PRTBOiBneEzwu7RquA7A716ITgUgOTNdvdNl1bT7ZjqovQpj9I1nqakbi
y3DxbuvVWK390zF6HYRmh9J35pcf9uKm86FCTmxal1QlEZPxrFwZI7k/mw8++cJUuXsgG1Np65ZX
r45Pe1Tl8o1nFY3zCrMae6a8Ao6fmrNmQjpZir/q9DcikDYW2RxRn5cDUybX7yx/eq+ZAOPAjsXm
VsbrMe75QGWGFY6fisSOHZ9sGnAycQRsmNHDeKyr8pcRg9ThC3VExfF1n4sAMXiBIPe7uaRDulSQ
HNnbtNI9jQCowJiAhtj/A90r0siv1iWHBJ6XLFiUd3TVXEjpZW2YRYbrmRe4WS4OSEEbUDAXgIxE
k15n3XUC89NmQTOTV90P8PQy1fcN8RSofp0PYJa7R5DfbD2HNFqVEnRddVRhdwhMnM/785s61jQ5
GZqpAKGYRetNZw6D5tQjj3TCa7fPQmdQZNdrgRNTGFMkhVO4RTeXvvMGzd7V+U7sEoBbWCmqVS0r
Zmi/NyQG87pvnzvhKUvLDtqRI/+2od4ii0qAJ+99ciZ8UQGQHqB4vO5dk+Hlx8G1BXvLeqMvm21r
DXGghPu0ETiWJ+960f0Kwh0Zh0n+7EvbFpwdsU25ZnD8c+7JLivHx/02kjSKhIw+UWklGF2qbMd6
lBy0Uopnbv+eDMKjCpNzpF2k/F4p5de1J4BEg2y7NM2N646UpnpdlwuvE4TzKwlqG1hXWY5wnvMD
mkOhkd51whFE/6Rxdiq+lLJ75DocT9vmVIV5U06XmezvNEPp3LeCgau9PUVG0Xsez46vG1IeZyc8
efDlPrIMU7EMLSSu8P2AP2Z3rZwlbdurUE8ZeYtsKJkjKvtN3phjSb9Bc/blKWeXfZ0+ld6IYTBp
+M5M/cugiW+wV8kc7GoTpJB+nIn+daOAoTg22QGGLwYji+78jbDJe1VaDxjA+2ILWbYT28v5xT3q
SXtRY+3/3Gps3pkq2JuVbtco0i0BjUEUZhVMcW2UzX5HKvopldn9f5uiXyZH3CAW77vreZSMCLJU
ZNWl3F2e5ZZrHxYTsThvvaHyS4jej6rvgRK9KHkdQGNIvHycxjvtlMQSuFlQwuQrareEIjd5RwIc
ORfDYhg5kSFT8lDM7hWtW5Nlaq9SLLqhtTUxVtuvDpgkcF/bmZpzHaaVosN3bfqqSkaGY1ksIWNS
oSZXClf5CURK+DPhsZTdXSMDsGi0sQPE+Gf/1uUoYdZ8cI7rZ+/AlJEjODjMFpY1l2w/MeD4A6Gf
KkTKoqlHMBP11xevk37H0KSOlFqXyTnLAucrYEHlSIzL9zd7BcJunvyeRBY61Y4+BIe4RpjB5BRm
CAVxd738gIgN2Taud425NyyjQx1K2vA4f0L4doJixZUxWqr5qt8gv6iDHlcuO9/dFRZIQjdHqCh3
B2il/aUr6GgwHLJYUkukCLII8iyNIoepczpNCDu9tccD9E0NV3v+Vb98B64sQYZtweb+0jTXtJvd
EHzO586vF1c8vkkctpmY/jrQ+Z4J6WSNjONHdjwXTunMjWqsmQX69lJ8VixOfZoCtXzxcy9q8BXA
fhaEhdLjO7oomNKGkiRrGQByQyOXKAhRlBAwOzrUScS0SOegWhww63qP557Sdb5kb7ElVcclLlfw
Kkx9nkex/yXR3NI5wFwrAIKWADt7i0LZijh4Q4j3vmhoCxOF4y4eomccZIGM1k/ETiO72z4rhDu1
lkc7MDFGVxBe/DLWaQdCSo63U2e3aMU9wK0h4pzrbZ2nUapP6tiaGbXhgII0sbFFtHt8WQJue/Zr
fiOaP7lH5FrznZysrGniUlgVES1/8p6zakkwBt8axNCM70ZrtkYpukxxKy2e+vWvBfmvoI37uXdk
2amculc1f5u1NWRYhdELSHYYbk8/2Vn2/I30DurLDHGCkr+zoAB6eBa9IBrO+hSyDeP6VWDktI1x
3eY6U+U/hCHt4PxDkfUF2uZZG27vInY5rsXEh7NwyF5zlyH2jkNQKDToROGQQJcBjcNerjL912mH
YisT7XcFVf9J9DVae4W+zQRrDTlzZ1IP6/xQGx5JKujsG8m2cMHSnEF669QLicJf7ZIeyQGJ7kT+
ROLy8Kt85OWD8cvUudrrcBqC7E0bUmvJpi/N579v/qEDpqrYttV2C9x66ubS+8yDrr8o+AMCQtis
emoaMSeB+whwlTb+xuKFV/B7cA0anMgJFSqsxcOK/QPmwublofyEReT4Dy7v674ciFKmVLuSv2BB
f3UIG6YZv6FeyXpC8IRNE1XEunuuEfkj9LmCzap1GBaMDE+CfZpp8GQ3fg1MpjIlxnyrWQoAZVf4
WbID7x5rrBfLbpBFxjj/1HFlYaxscKvKAkjmSNCBwuDYa4L1dWk6h+/GMbZUYepmuDH0xbf3Tsx6
lAy7d0lYVmVvRNbHYehCDZadlvGgv4Aq0IxeKo3Pvy4lQQVeRNZcjksjqRYGwemnnoumOn3KTd0s
K3tY24vinGSGo1uGhmNVpjN/6DFwdbE20Kkm2u/91/BIwoLqSEm0o0hgzHviC+QkRHhsHVq861Rx
3oKf2F/bHC7IpA6oFtD8ySVcKRhTQvnCao2nAwY2Pe9bNfSilMhM/JrNIJv41GrZjo9E9B50CyAX
6ReJdu2PQmFeeQF1Ei7ZQbCWTlxH6K+CacOrf4EKHNAZXCydKU9yJUhqPNfvzqD2iwZGRKzj6sZp
fYbM/pRXeLaJKfSXpA9PXz2gQkUvOQGT/2dqWqwKOI8x1dCnGDk6HyGO93ppM2Y8xPyEsd+D+C6K
gU75TFh/SOlIRhGF/DHK8JkUaaC7ND5nGSI8/CazYHHZlCBmG6Rri58bYtcXw3330qKm+cXvaEDb
pdupz5eIqP89Y6fM9ayGoTgVSZgQgC2+/eYC6GUabj+iKaA6Zljxj0ey1A3PE5bf1Chjz2GHdPUL
7Wy9xvUoYi7s6MKxkRzW8IwJHj93ifSQDyU5VF28wRez9Z58tfNVjf2YeQ3LO9BWxzjI8jm7bpVp
By99BF/1YxedT6qPGhaN6lt8ru/CHDaDPkRhSQNhr9WeF/NbYs61JP48aW5wIBTxeu1D5+F/Rilf
apwMKK7zWYSAkFnA28sgPbHXM3EYSM8rbKLvpCgQsOVcon53tkpBoiF4+iXywpFkU35UgVkhGLsG
S/quc2YJrBp7NpTh36zsuyTtwijFnnOppkbvTZu4z3YG0KDlf/ahUDTK5PEzBL9t93hSdCRb9Q/t
k7t0li4MA76zM4xgVl2SMFEudFs2u1G5EZvRjLXsaOYjWEfVojnE1tfD6JVVsOYQhGWZ+FRX41DY
mlsdJdOg3/xMNAzVcXijNdNoalUDKVxfrdtBTUVlNXPj/xmzZcG77bmqUrzpmY7U47ON8UDnct5C
TGDSgk9AFTz+keO7Xq9RysHRrwxz2pL2/19HlSj1hTuCImWt0rC//itOXjWCdBrWIwBnQnu5fFuY
4wLIyrGCuiIp7YgV+VE9jlOMYluzgxIUu6uNNEHO5OcYWHtbcYekjDS9RBYLrDfJOD6OxxFWv4zA
Dz8tGj4+o97iy8aLgcNq8OusAPHrdzLdei91h++mZSd/U1RCiXyNWvOCYRlcm/VLKF2pnd+T5quD
PAMixI/iJjfdrrY7IQ7dn7nIXYaxgDA8ZrKvdOPomcTR3xFLrCuqnXSjlhmvid6EFvyGVwv5yYTS
eqDSQizED05J0YySVVqmj5Eo++H8sustnThukWZkB85eEmKuIpESqx9wdYMydDZrRXou60LLA1pS
vlX42Pgj/u3d6RKfw5v7OVsQbNXGmOH7eOR59a9kQ8USSghfRPdwE4ZAyDMWD/MwKwuINEnY3Xan
OyHe5M4QWtpC/FTNZXaYL4MdT4ot+mMwSqeLYs7A77iuHMxqqjWtqedl+x2FCbVD3KSqnawyJzOd
nr9WvqQivhLH5W1uzqRpOhyM9Cr26Y8LyaEWURQAH2hXbNNBm/8HaXJe4o7KYE82yr8jwENH16XX
AQhrL5y0/At27EhqF6r8IaalB5Fh20HAJko79S1l7N76B8e4Z6XLAQXxP61fnH7kuteaDozvUfUZ
1k54X5asVrT1wQSv8d0XVzJSr3U3NSeUK7JmiCdDYyMTD/vQ2Pyoanedlp6rs9C+WC68KiWYJAzT
xSDL/NjRpLUn6RIa9jov75EI/Vhq+5ES+UQwykNtMuTf7WDjgu1b+XwLyoTitEtMaemtuXmJA840
+uKGPfUNKPT4qeEZqeTgHaMYT/xCYnTHMeZR5OA487EzjsMRipMLSamgSwoHxXYZ20utVWKZy6c8
YxVtUisuAYZJOI4ditM/DsLH6aqEyME9ch69r0zlwyryt3Gfe+bQyuWhHPQIt7KYQ2PaAoAPioWZ
w+4FvFthrA5cNdjwwYTFxrASk0NNrk7oEVaz4KW5s0TWUaqRoOx6Y+hI8HRvzB0gLxCLY8JftWoi
aj27HKTmQJJiD/46tkxSmLwKryTuEjriKtrouamEx7nRffTEqaHbOIR0TXHO7VZJbsIwGGi1Gpud
PElUQ0XK2J/Pp/X3Cd4XUKXBzZqUqOkQTazwxz2/hMK+lwL2rvJAUllAdf72YKURyS6km4ZHktF1
RPR55yR1ppZXkyozXJYi0YJtqR5y9qtZvfQHiJW/TQE3hVHcW6d/O75o6tHz0FgRDS0RzIaYdnzr
NmoB1dS2TIgrn8X/B16YTM3ps/FAdz9bmKFKc6h7SZIT7abMM2ABICtnA3BPAoo/JPOLEaNVXGtd
lVUKghSCjgPwqXBAU1EkhpJlOvUH7VLn9Zkh+b3wnj5OnatTuNluiuysq0SINPMNUfq1MnsLKXwK
CBHScVgsFCiMO9bTVXR+Q+ahs8ExQlbAA3wzB0bUqq/KCWso15qslhY9dJwgIUr/wwU/G5Og9H8X
3W/3erLpI3o07GsE8rhUS9KTr+UG6xSmyfBlVLIWa0zlD1x0ZIOMH7MgIHo9PwQKAajXQDYN+Szv
zzwHpmtf+0wDIbV/ZBN0RcoNeQr8cd0kyZYaaJ9Ut3Dua4l2OXnUciOLaAzP+ojBet5xTvsLAiyG
HiUFAZY4fb4I/AyUDNG8hPyINH/ZzQvNcfeoStRrie78GKIOsRjd6S2SDAB5ackvX9Et5FDQkMtC
6deHrdSDievsvfnlkDQos6el8JpSNlY6YaClhk73u2jLVxUyoMmTJRYZrSGDAYWJ9VHg8JEweaIH
6fS7BqIRLOuMnKQnGB8YzHd0GxjdW11LetThzGcY3upJNXVb0Z5tJdv7/A5pYD6pQcuxCLghBE4l
7HXuYxzeGWMPxOBkKUyjGZBbDPPyEJhLL1rI/OiaSshhk3UWD5IlFQECQWiWgWoVhhnpqleK1q8a
kXtGraYX8dTSgTe19mtkSEEbLTaubcARZhz7ji97afxBqx6jSpajnjouvfvdh8DqvOFd8LKC7rc0
km9DSd8SDcaylpOlSL+u4B/0MzvuU72z0OcYYOdoFzAajyS/C+xB+BlNJ0g7FO6oxgsdD3QxEaLt
6GeDwnNuzfTKG5dkgRce9CUsqcn1xAiXbf9yw7oVj3xv2WnxqUoi22MRx6cQNBltIf/xBhSdp9bb
gOCTop4xiVsBgJbWHwbn2fGLAsHoid6P0pEdbgbsERy6LAysrmbl4p9rOlpqrGL18hPBa9IuPfC3
c0jsThwhIQUshS+GI9Cxl8fPAYtXgyIouN/bFu9eGyIA58+SSvAtWtMedyrZQRGA7YVX2m3tG5ts
ZOKa8PpEJhqnCZSga2vVmcBEUMI7Mg3HCOlrpGWd2YPvBh+Jwlj+FAPC/9xFZ3D4RigMpVWerdyL
jQvNRYptY5sW+BSOF44ivzFpNMPlQUFuDciViDG6vYU/9uF76OOgyJYg30Qg3s9AfBpb5Mvl3N0B
vRpqHT3qjupnlRrH1lSYT1nyKMu0hRyOSxnEHNrA/fyW7mcX/DeZjxr2vvgRx2FY5f9fs2Ws/2S6
AUJ9mWTcaOkGs5qvO/dKePzNmygcrCW4nZMFvCp5/VJPU3/N4YtzobJL5lJ7QbeEgQ90W9UyhMtw
x8vwpVjV1ofDhnc+LM38WQTwmOfwLAs5RkLLR7RJq0IJzCS+DDTMPI7qXBholbOk24KRW3K7Aum6
hiEqJVWBjOO1muaYfCtdDD09rM3U0TUHXEYz8ZkOmgCdfrHYXQFNhwiI847pw7WqMpmfeZo67OUe
OtInwy6m4+9kRYVOepEPVlgWq1CtBXW4ZwHx5+OHKzuT5bgnEcTjYEHQZ1b4jH3RIMcmou1DDs0u
xr+a9bMZLTsf8SYVig6B2SL1K9EZhRnU2uHfAfNQMVlhOYm6YETZJKOiyjahTORoZdfW+oaMyrEj
7/r4pIzgBZ0w54LKhashsCRC2203uOzpvsGj9zLSqiPd4MR2WH0J9e12WxEhKBlfVGe0Fe3H3S+v
255yuC1kH8zIb9hkQj+OVgLeQoMnJIc0kFoNmIBvlmmmAM3r5/H4ji/Nf/U3lLlSfKAOVYHVM6Ni
PHOoV0R9irs9G0re3ZRgBgtc0o6/BOpjGKEjYB89xfRRx4VR9nSvPLoRnkbeoEkHmNMT0YBMxE98
8nbYUOI73hOIpe0ZeiezWkfQXoB8D+uw4fTAwzKT3d+FcSlDjChSk0tn5izZNLFHUrb0YD0pPQav
wNgv7UGxjzbx7njVnPmivhOpa56ODvIuU7GK9JITQjMExotByjqaPZf2lajEsRS+UfjD35NUjb6B
BZKiWk20kE0VI8ps7/nW5aE67E17N0hOK2hByW+FHsKB4ylbH+XLU/ZTCTLmOkKesVel+jH9BVXn
ZdTVOZU9iv6PpkfNHJOh4/kl+VR/wMqmKy9kjFO6VagX3zLbrhR/r6TULChKUplsky6A66tSeobz
BdMXqtPPstOfSdSqjthtRzhGms3ir5zXYgoEr8Ii0sr4ayapAicyt7faTqLYPqC9E+OFveEtxY7n
YH1tYxYcQRJWTnhQmLdfmVbnB2mRz6KCtGnMkRv6afloQyWz3IhHhQdoGukLn+q27/gLzh5qrY09
mVhVdKMaC71zMHc32//9GpbVWpMV5m444QoxBvSFS239nodFHfmsyxhLRnVS0d8+nEc8MdWJo9Mv
FClhBMBP3dNXAfSyKTwhitQnPfdyz65mPPZI9vU2Fhmvp/F38pDjbnRmG+gsJiFoCt34bDqQj6F4
DtRz1hxefpJbZNtkfnYe+Quf7TuHeQL8kV7+WY0rCY302C8tlMbmnyEq7mgQ2FNZ3Al2T17XbZ9D
+tFwg+NV0xUQOKeEUsHXuNf4FurlckkpsjTh/aIHuaM7pjiPwRQ5/qv2VD4BIR/6zocp7fsVWPkf
SpWBYGHQLAp391QyOO1x/9qvXdGa3T3yxpi2qwqSuiCYTQ+iF2Tc9AI0cOcuXpD8yz0H2g7t24Lf
NjUyHhJLaeoXzKB97YCQFg8U1j+PmRZT6eC8zcY69jyIoxk+A9xSCt7eFMlcAVinwS1Cv/sUqGYf
5fleN0SKj4jdPXdX1tLjlAqPtkVohAjC2Espre3dVzuoJPIJFqckBC5RbOH5J79xWsEYEIc60g+a
ie9pvCFTaEhSx/dv+qN7kTfInstvsPDZMXN3fgPylZOwDqI3FajKrBBfJbsKIqBx8m7cPXZFx/vR
zOiIYUU/Fi/iKA33yerk1T9heR2TEcT91rmxCWMTCabyupJeeqdRC+f8N6jLEPuA78FvJjyhcVHq
q1Z3doGelO6efWUD/g4U77YlMJKFB5bcsy//4r9ew+AYg30PCv0vjVaIvC0fikWzIkFhwMYeoCyn
WbCyxUkB5sH1oULWD2F7KnCZsLOD3P0aFCw+ehux3xSfnZqYlfYzm7t8kgBd99Rba+4jicEv3AOo
zPuA7P7YozRYCzazKpU/rFJ6UvqVq8ym3yJElKT2NJyPRx/Ld9bR4CUj/cSyxuUqVTK8A202z75c
f5eeom0bpHMNMRY/lihjzwBjegZY95krZyg8TOFWB7gxqQwBJaYRFzcaXEoXFVog37fbKqRSuM/o
0Yzg6N4gijIya0icURibwMRD2cf03kZLMj8wLswrJYY9WUXWMI24Uc7qSLhe102hCGrF9aJ7xWmO
utEC0jMJB7AdDCmB/GtGvjjNnc9N6VmxDDJAtQqAOBxmH87Fw6TmG3eaMfBlD8P+wGWo5oPX8uoe
ehbmhxdoM36lS/ZWlhv0JMZ955TmE0hybEDi2ydAh1+OeQZXSE0vs3WvIDmCA88XM1W0H+y8iX7t
bg/orZ95VH6sxUdcAICDjXi8ftAoTbsSRJDF3CrbT9/GQJETGyhqLIwuZZKHMR5DT60bLOYl5Zww
VKnjxm/Wilkne0SvmcvgwtoKWVJAuAQpsOUj2+Uo6LB/LK8b7oURyYMurjEsmwzPQ6AezN7dqmhv
CQLjd+rZkruMgVOufcrinVHMLGkIumTlQMODcG49IUH5ggipOLaw/ZgDmfUdhAE9Q4oxxI/SISyq
tn/p0RZgE/K8r8/T4QODputuSlGqtN/d2nmm6fgO149TAmkaPq6Z5jbMi4MKA1Opdmcsji5X/tZp
RG6b+V6Mq+t6ywCZPUfO5y2kf6idE+d9VvvrDtlJ92/Z4XgO9EMFRKFCwMHaEnBq9ZGh3CNeyk8j
+TKixvJcIQdKiYeUTWGR/tPwVV0L2br6szusS/teA/pXOAWdYQR060oBMCSk3PrabR1Iar3Xku0T
Of5pYu12eECrYLfmeTg8dnou+m8MCzJ5PbQ2Dqmi2WoNBQhg7AyZH67uKFvddRmGuvxUos4KIwg4
A5wLdKDkYaHhQP57gC/uMQ4kKdRCIMkn46JkmLV7UCzgQ7tYZACY2lwxtyV5uOtDVInocPyF7Y+e
kLzfm2wiWXKQywBZTmY/XMHIDYUJrydr+qg+hIXOFwRdeirXsb4oHPVwpeLfybEViFK5Ab8uaG6d
9PTePddJVLYUTYxNEsD8Jz2a0GYSjJ5TTy2a4YREkzPtbvlD1e/pyMm3TECk8qS50/I/T8SA8xU7
pzByKQsE7+FyoQMPgTZUXtBal0Xv2SD/Wl6xqjEXT1r20JFtJinZifPTVx8fnbAop9TO9uvT5UBl
I4E49Xx+NjphT7zBaHGOtBLxpgl546UvQDcQfbdN2Yq1hmubuZ1nW/qLQ6sqVZeMFv7GOuGKDhnQ
p+3nlfziIJCBAxp8SmwdaW4AM9qtrO0b9MpzLiSQ32Xbs/W2mcajh8l0JLHDnMsCqfawU5k6uCog
3oHO1F+/mStQ/jlXVUmxZ8eT5bPir3Ufdv4QuM0I/DpAVK3fr+79Ehc6tE3TpJG+KVHBUsf3QC7z
hcJIwHdUPxDrcM16uviq9rikoJGWu8FRA90baiUkAA+fF8iQC+cC52ObjnSZ/mTCZetW9vLtND6x
lWFSPU8KSZeZl02FJj0NyFx1T6/jS4Msbb5Y0aaOPxMaWu+E/X8aNpBFjSddXE3EwW1XfuZwolAN
SIc+F4mf1CWNGBvsJl6Q7L03WI+eSWdenOcLfu4OAATnePjwwcqAEKpZzvk89MbyL9tSbaqaJTmf
jGAzOP1v0ihWpu9nE3Z6ngwBaJvrfPZkrp74CAtDUAt7bs0SX0Tqqfzl8avtagp/TblRQzL8BQfE
qOeB9Z8AA4qTO249phuLC6FWxBywqrqXu+ayOQYi5Ir4k/Ai/j+wAIfIuhyaUtrZ1ihmtyh6OVqO
yw1F1aDqHti1SAzg6Nfcua+njlA49m4g6pMtaV/TFgV08bMCki+jOuM02PChLYAaza+SNqeibTYD
FJOvoFVk+MNtiCReduUO1ZhbeszawJkW8En9mAuRNDpNj41HegPJNQ6shhg6cvUvrH+vpJK3CRww
8CvZ4DNV6TszQKA1ee2nU9ZNQXN7vXxBfUVt1D9IwiKtLX8wzDB7T2ictk2QWTni6MnFP7buSSGC
stGHdyNKUjVK9vymOLVvD07nvmWRkdPol6Sp5jE3zgIAsKVHeafra9ZbOFkh7UlioR5bwHIo51iv
5krDOFX37oFdp/zoholhf7xEZQCV227CpdozHfxmBmSatg6x7Ag5OJaUwcu2qI8tmJx2gKbNbciH
lZQ3utSrch9TOo8A+Vb4RM5qbfWEewXrqTeikYJe1DYxx/3iB02BIaNcF5xzJvkxS9d1yf/DBDI0
JCGslEdcugNnr+6gKpMrwtak65TFOQGl3zktonOCfFLLnHmA+wUtG9hr0rlsm+Y1DIrnuc8JbCGO
z4Ys/kS/r8yZD9aAIUWiomt8+1jv8KQlGWzREjwUis0/QRqyx1RibrKXv4EkhVjtB4sgqlgXfn99
83vjEgTK/s44Iqany64/+24EeNCmmR5qC2CIwFSD2LlE27+SG0643Sa3sC79zaMSm0WkLxcGw2DV
yp6oXm5sXGpXDxc+Iq8dBmJ+jKTNTn6jHXTiRHFYzvEPAuiF7bcj/tiA+e5VWzvw6QyTc30EOnyQ
3XVy6alpnlJHTMC1H3dpoiwuJWMsNOgPnwgcIEt0Q0t0EU0vX8SvsWSl70lYIowLFoMwNwwbMYAZ
V8OJ0bgERudsf7YR9+I1aGg+SQ0yPPY9FUDn3EMGo3OSArrZEdhQonxTsE+5ComUlxCOSdLEWj7j
YZHm9+DM4KJ44LQkGW4FYMHwwyj+QEbX/HFzI7y0I2Adln8sppbUuWL6kHw26SEerDa+yX/EKojH
Iw+teD38zVp6obZDwaR0cotTLF03V7Br2lbh23jLJQmbpqp1llN4EB+jcVhvckZK11qE0z5Pi9r6
4qvZ8HFkDghxfWVQpmlfUy8b9fLjmP7W6mtmvEnxfjFxLPWSnG4D4zVmBff1t4OLzySDDuCfPiRc
pNi+dPTw1H8nWb3rOPt6oUyqiLsOj7cR3hNbKHUQWGvZgmWi2pWUTWeheoU18MjEs1hDAQ5Hi8UR
cFJrnpaDTtTilakC+GqXuSyUvyCgRS4FcPK4KOukySIyPFjaNZz3zVUKdASPdyAux//d41f/iVYF
aVDfJOqSgB6Eq7cDK2PYq4wrnMpQodaQk3ZH1Iq/lu5Jkvx/pqPMiyJQGpETsY9MHXqt8p6qdjCR
28sX77NEwRgxbMr8Quxc/7N0qgcTA4EVckvgpV2uWp9VSyd7+Ktnw+AFGzqXwYQ4I2ucZgjRiBx6
QStliKxqwYvLdnWs+WCikaSdaYpjn87bU5V2TOEN45rIECcsRA9WDjgMUi3fdGQYFy0pU8Uewlof
yp1lw38jyh/y3JuOcYrT/ueVTwnWstWD8/Tv62ArvXLagd2HZdmXLkmme02qOHp6q6JsT/DSXkb+
b7ITMi/SgnDabZqnTsYX/CDAtpSfiEnaNHRwbs+wn2LCf8Ym60VI+7Q4J6M615fFAzsH/oLC01mb
Y++03lu+l3ExnqDsmbkFSRMGFVc4UJOc+8QLQITsYIuKh1oOReasRz5LITIVtLMgh3nSYALeq48n
sHr3MgFC2WfTA/hT/XLokUYoOC8NIdVBKeYBNRemH2f6j/H42bOhB5CcveTpYCR57uelsquVlCBy
6hQ9u0oHpZSvkhB4NdnJNTGr0jlI31roebd2St4nGPVW0x+ES4/L/y/2gZAFI7QCKrn1D0uXK5O6
ZML/lQ1fe+vSPdbOiFfsU6m+TeYkZ55tY7pkwENCm3LJaCyfmqiDFxjUm8fkDlacGwCQOVuvUROn
vnZWJZrb8fxwYCJjBS54DJGLIRhv72ks87WaQgdsOjfKRFK8uZCT7J/FxD54bpU1s64zBS71lk9f
y+CMfdXKShd7U210Z83wELMYq2OFaRZGvKGRg4eaLz52PAiCN7sHGXo25y4gid3aapYHbYzbUouU
L4nFz+tGYZlnQpWI3H5mxzGjf4dY8OhERguN4xCehInCtLT9j5/JEiePC5GtM4rN1vDol/47BtYZ
lCnGZKJdATievYhR5TXbJXafzWNxUG3esXH3fXASkHJG2P+Vh+tsz2l0RQ6/7dWZ7DU/HYu0koia
JpisfxkWERjnMmccq3ceXSh+ShF8KrGNphGS1ppBdpRhj4i9RmfJF3Kyw7iuxaecx1pBhPyMPH26
vbrd0RjqVTCoSH1glx+4HpZZt8Unaf7+6PcCst5bSFvfaP5qiwedtNnmwi12vDL7AWr7FfzmOM/h
oTAqa1t97FZXfWi3uOoO1pd2tN9yHy9uUvzTslSkIMa8gTIas9lpAyw7F6SduXkQUB98QMvi+71r
lS3Fv35RNSi3qMzcfYUE25HNPFvC2g8i021r9kuRKGTv58ClRqG3tyjOW1XLbRU0zGOACt2RB+0K
4eE/NaKKLPWrTAnw3zy/k2FwGp4VZQ363gpB4sLNKF30L/pQZ8cmaYBQF4x0KNAsQmKQ/AVUQAgm
VsaWit7WawixicrIi5KFgWlP3jVPaRXDSlG537ObsxovNSsEVDAlmWuAtY+T8YO33unR4B+Rwz3Y
L2BaNToxtgUmTSClUOOBkul68N6I+M4GejywE4G3nuexAzSncZaoDdJHKZAzgQ3fHxoWAsszzxib
HWJ6F+TdcyS+k4vWBn3/GtKug8eWUFy2agSSbCX+jADNJdxfsTumj8w1HlPOy399x6+51EZ2eiHs
ycQfDQUh1Q3dG7QaiXbhMsU3g1RCf/4NzcnR/foJGAHf0fa7anKovPqgkE+E0YsNJWLQOT5rz984
ZWhD/vIc4i3EtOY6M/HQHzvqrgUdabeNzzEKxkSwvrYWJLHzczfsdDcKfsKpBSORQxzt2X1FcogI
4bjjqeMVAPZmubSac/JaKJ3tCiJGgSssbSh0B724n6sU8jsr2ZJNvy888NXDCzbJGvCzndH1ED7j
y+i+nMrqHXkuEi6FDNOENggyYiW1/WKKSlhodDI0VT4++eBgZc5QqjJ316qNSwc9O0doi5EOMTXp
W1wvU48e2aOSRo8Mmg6/drFh41ly2tAAOMi6XOADKFvaf+cC7QxkDsA2VR1pHDjXHn5LDkVPNe/b
jgx1A11D7U9cJ7r+4ywBymUZJWtGIMNRujWEyLFagkcAOeCoSMl7rgQPUN1uWgi7RwR1hpykQ0Cy
AZvZuMSfcr2YwDd+7ilCQvGTjoW49e10qVtRFHmikreXdh/dtrBIhW+tuvcXhdymrrcL6kSiaL4b
3nBMiVxvUpF2WS84Z98J02uQC9l4MzdzkDAnFonms2/8o0/S/X+1aDF3uzRCXzswFENyBMyucg8G
Qq/3QFRvn7spr4LfudXgulOX8S+tUAYOG6HgRDgqcSTOAjxmt72v03QPbxvlogbsC6M/s7alLe7e
+PKAJKVrazPzZVw0TUrgcgfW6rr4wUtFJz5M+hfvKAK0NlDi1qGF2JJCcVsPvO1vrrtiMlP7Cs4t
Wrrmi54twBsKzacJPDpHX0AaxMcYFfK3U4hy9XIrzO+/ZyHVGC6GpAYfJLDy/Cvdohu3D06CStjC
46KnE/cckGpFFbHuWT0CttIi0hE45hgThjrE7459tlsVk4pxafcl3ksWYxnLVdGKeVFwxl43PRH3
NR4QQ8YorEEpCg4U+SKdmezXegScddpBmYTMCDi+ZdJ1Y3W/agx6twJGBXMRECJoxtDmvhcliyRr
ZPe5XhVWj2WDr2DXQxLik0Knozj0KY4QvQ1C169KXjmqZTWm8qcChmhihorGQFA28TpDouwpIlqI
2cSJn0m7sKEEmQql/aAtpCEzefXDl79JAxH0wOUwkKHbLkSI3JZRe6GrvRfQm0ScJxC3lNawk2I2
HRaxUdah3mLQ7NtCvqz1JgdM0ukeljPP+nYJEv7zg3pkaNRFxi5ElvO5G4pS2YMtjV0s0xvboFxt
jQIVfM30RE4gQZDlE3G7CvApD1O/fqDByfX+QPQa3A4Lu6xlI5QZA3JN0kD88+Pe0Hfu7hpFb5n4
PvVhkGUfm6P75d4jj0zcwpQMGgSs8CK8smKJgQIO3kforMtrpCVlscy4nJKSrVhPNpb2D/NSRm5d
PNSefPFtpct8XV5c6skR1cfntOtu5z+8FFPTIidg+8Yi73sRXxHkMOG+vtHwHUZf+UFusJFgdyKA
841ovGCTt8dm0PDFSba/FQG/HzzY153FIkq8FtXMDNMEwcibWY/PqKdo+kc6DVLD1WHuFZ6zztve
FAcu4Jxg24x1kroMgQ4vfcxVRgVODVM/NhBYb/1DGEMzS1UTaRZC1Ys7Uv6CB1NM7pYldIA9BLfw
XOtrVKkpJVH/jF5IkeH7/QsLyhVLbyo5dP6+3KPSccF+2PW7CJoachK9SDatY4XlTfLAJbP8Cz4K
b5IM8WLteGG03kyWe9KPcuLKaphHpTzkn0h5Q20KLPkzIOgx7A1wrOc9ubGRAD63fCnuMAdx5DOy
Sblu3SRT7zeZEfiaLybOSOHm1y2rYXnqYpqJxr4I0DXEd+ZzoaNt5NTyda9z/eLxIMERsnSCqgRi
BjTJ7tBnLz9uNYmpnratSSfINKWdjwTbWrhau9BGdisDY1lXBlQr5EufOg6Q2G4yEy+MoxH+3DBZ
rFU/kXiSgk/zgT0eLK9fvBhz/VCW6C4bexl3jNiqpxERsNHYS6V3cjryOx2AX3WZ0Fx94SQHXQs9
4rpVMxfTo4T/+ifagWr/kv/k3+pvOAKxtrVK61hdxt3gmAzH0NYXD8eeDSbLai6CULFmZvbrHY41
MyVYqdix4hUGbRH6AX7desWfRUVhb8zZJzjA++qQOgU57ha2PgAhdIJpskgzxBHy2sQ9OPB++POq
MbUQaO81pfFWKVcpLZuzhA0BMdZ33WI8Gh1GzV3rLKRdUJdoYlL5HDj4GXBZ2vWhflSfzUlJdW2m
uDGvr57ykatbvlcRUp1twCAx/u/2DPm1klv6566XHjp7tKQt4BUqdNrc7kfTWjp6Cwz02XW3oLmK
GnJvBwq4XSN2neKALR+Qwa+jigZcErYCtTFyeLse+vSEX2fsvHOdZ38pnW2JJnynxVCcUPBDjreW
DOSUPZY3r8FYUCe+5PTYa7m7cIoQwW08Yz0uFnYU9Mc90cRQGrDSNH5vsFvB6ekW8C7I5IGzfWv4
kE45etl70fJ0V+vjoJ447L4lR03InX15FhQpxvaB7STH5J4YEBMYtrEaxGssS58FhcaJW4DrDSJ1
joKyU9SNNGKtyiZKeLUXi1ar5OCDXwx6Wg5wsl6OhohwpjUHfROylrLRqpzU9MrPCI2jgqAkmohl
jCbR5BidW500IRy7ocKWs27vMVT4KkLMcqir3PClEvO5YOSHCF4QeaxUbpLXmpdHZNb7tlXj/w6d
/kXb1gxKuDmJ1fzWKPjy1xTnm73/SPR+RnTd8zPeuqn7Wp3gSXiFH2AtV8HamOCCXxOxRU+ZgsYt
kQ/a6nFW4kvOJ2fTxIVschzixV/B9ncDbw6JluX/fPWjtB+/zTDkNvye3k2a2Zz4txUOo/AA8fHn
nABfHJQ8gjbJk5NQPxAg0ViJJYXwAPRoJzNjQHj+OQYosTaIYzOPtqgkEi6zmPTGr20en+9xgE+/
tIdINuH8DuBYJNGCNbxHmXHQm3rATCX+FURRbbUzmakhRwUXwoGnfhkRBm8fV+8RH39YspwaZtIM
Fg+u4rsUGBDou/pFJbHcRJM1XTXiuufp9Fc4dXMttXu6oWjw5ZsMEjCtVRFcz0AEfmNx7U6vuR0K
n1MltOM8nO4C/GGzmZund5UKezlDyUk1IklLWG16F0LFFeAdQ4lrFHvN4nz6TYtVq3UksEbz6blh
kxPUHK7um6QZJsZEdsRGgGmahdqCPJeJzW7j3NKSz/MUzXTdHNxuA1eB4lmMtwQ7BrCM6K4BlxXu
SMQOMpMnA3+5nO7syh0JheXeZxSbqeujZESgfam2jtk9yE+/3X0vZ2Wkdh3u+Eok6Nbi3mL29oRF
MKshzJ6uGlCG/2mFXgpDJCpy35WiNJ4OHAAkMb/LVc24m43tYEDjBGVqWn70DYRnqE4w/dJx392X
X8atLOZJ21yZOOjM7T0GFAxkYI2+KTPF/KZ28ZInPPJKyeNkJNYTEaWisdN9U7q/54MKTao4qfE7
5WQbIL87gn2LufBObHlcYFsIx9Uy5vl0qtqA2oiejBD/ZduQrjTl7Ig3wcyg8pSG7Pb2FIQ9mMYN
HppH2Uwz/AJHqN8NlFLLNOL8r64Zspfbp4ak5OaOi0h1ZDFRZYpZsY725msHp48fSlpwcVi9ee+G
pl+4vDsFKE3mcRoQvrizawlkbuVxSA3qVLGH1Pltkh/zcJRGsElpZEpfKNF3xg0vYdzWAT06SUYO
/N+7poCDKZCuhTGI+DGhswIpo01zm8WQHXcA2TmwqaOV8fc/iTAx07U0V/57ARwN4wvZbqWAc6UR
xp8IiaqC01Z8gnw1QF1A5YEzLLeXsVGzEZ6Ba1nVAVUBxxcYLllcCnW2rrLWEcazWe08GiFh9zIx
rr497kHiXy+e2pkWTX2veMp9XORmJusdUF+KKjNud+vi4msd5ZzflUXkzIXELvjen7XbzsId0QWt
m+rEaOvmNWxvku5gaDOKcYP3Y4hEFeHoI1+KFL2iDOXPwTXG5enjOnKykCy3aabsMjF2stYqC61R
VqJlFMBBPcIE91GlPUvyen4OeZvuRE6+40znkeo1DbTcpZ08mZ6WQERMv4EN7UjiG7oiufpDDBPk
3cMLkTHvuOOM/sIJ+UU3w4XBAmnX7Xtg+X8GULwbW9HN+CK52qzRsIb5/cQM1ZR+/GVihW28JpK0
PtRhxUXzecnBxH2mdpmI8j9olzRx5VlQv/7qf/6OX5VbK0MsQW1A15eqT73SeQ4HRcO89FalYo1M
nHt7EBYfK3gEYAE3dMLG81a4I6Snz8DJ1eKk/xe/lpP9l95SAxcMkbWXDwzjTkYsY4Huf++0FVp9
9Qu3xE6iBdqy2qfz3HEsBq7ElHCK0U3Fn+4ZohbaUuoKd5YBy0MhuzHj7aiYvSk3qxy1brVwJ0ar
jpGBoXM7R68dCLjNRQ01dcpt5+14bzzPYsOfPRy0XuhxCZxc01cWwioEzkomzKyvXW1OMDzbbIGX
kJ4tng/73Gi0NZe4s16hXdIfWbEZkGfjODdv1PfVITUYGWQIrsr1riIWYcpotO/NFpBXgzYlMUy9
AikD2Jo0wtgG6yVBy63Q0IMCUpGOimu1mtLYVM7XBymwjgz+ecgY3/LVLgcWT8ZuBZNnIZxPMey/
puDI4GK4BddloS6OPEx0HJCZeR/jaIfyyG7Q/PbctGtqUy1TK0xijYbaztr8fW+1LunwQzeMMT3R
3oGBmgXBSeX2LNWI45hDLqzIniJrqZjGsdvS9qSZXu9ixysmwz4/x61ieW3YG6NsY8KELDVRoqFu
CwJh4TKZqySPcqJr7WCURXEXqHblefwm4Hq1VE/psR0Moec2EswWS3vG+H54qhMh7zmTqtuk8Ran
R5A6l/DLk4xWli+3uADMhcGBFC5VxpwUiGZbkBmygswTcEKCRz2faT5ur6k6X+gYZJGg9VlPeu85
wGuKiq3xZHay5+oNEvv7tyNMO/xEbq3GKdXw4Lpq8x4uIBu3LG47cF/um2ZtA49HPn+hvjBgPW7l
N3ZIOqNFpaUi2BvTP9pe+uh9cdTT1ry7KmU+gOaoDmeT8sv3N1suOExnu8CvETAkDzBZNF+Sm485
KOreedfTCdIQ7/V43aSVbEHO9XpMvy+KsS0mvv0BD8Vum47ginT8t2UeWW+N8tASLjbTT8rDT7zI
b8wW2IyjuJF7ZQh0uT8hlCHPRmRDKu58Vysky+xJMwVFP4FlrJCjEVkWybULkjuoxD8GN+XdHowO
MsljH1owD9iYRifQ5TU38P7TllXd07re8aHXqm8pzerwyPXPHS19OI1SrmPwzqO+BYp1CkZVNEmD
qdwJ45l0VfcSMTTACxk2tHtYOYXJ7C9Dbcrws41mN7D8v0jrzaCj+NPlNb/qvl35BDHAoT2H7QoZ
OxpA2CGFNUQqWIkwPqVio0UgOmxx2Ca/oK7g1Y56OWaWTgf4t8MWghwvUBbSjvmcbZUlRfAuX7JN
ZSkXtZf2scKvw1p5F1jdtCeDWXDUE/4vUBzsjfUPfAM2yKoG+DPev+Z1gmswQxSiHvWOAXHuETYm
WYFjeMuP35cmrctG0Dc+tdbGUVkt1PXC93O7c7C6VCIV0rPChj8IpK4ga1CBJwr0xJaMtb3BXQ1F
xhlAvilmXlnfxdl3AlFxWecM0FFkhmLNGLfu/aTCyJdXbWURTU/tKOO4m/Ey2JlzndzhhYosAfUZ
kqTpztubHq4snBVGvorcb82izol+lhHVy7tewwSYXygK0NT6EeBqZwzv2gapNZz2kDj3QKEM5kd1
S2Gc7YJdUTEQFSvlGyiSPVU3AisfaXZW0CZdPZbCyDv+P2BJ9RYEZh0QQYnQ0qZmiSbpzSIoELvL
vwOUgUdtTNklBzY/G2xDuzFa7RKhn1Bbf2Rx5KY52DJyAmaqi/RP/KJqriVaGciuRD70XzIYUnaA
dY/WPbqKqs4rdhVY4evdpRLYaUzzrxc696FGUczTFLJOV9XQhGroPRMQCIPVkQ1hrrjtgFoErp8T
ql//d9kwx0oLiPKor/hac52IkuhQKZzLyFsswZwBpg7KaL2hQ8E7Hr3Rn2HWRydr+oPoPXSE8q0n
tlske2cU6ZjiMNvNetYrRyQlkZQBmqrKAWAr3uXIBhuGqQmSxzeqYyidBSuN8RSZMOH4tpKYwL2K
LybkVy+URGQVtThD/AB9W65nn0TYvhBYeuUseJnrlSlZDNT0UtAVEtHYqK4eZbFklQ9rTbFB3LQY
KIxMrfRji1lzDBlbx8vWPmc+a1nalxMj4dezxWwaPl67KA4wl7oRbU+Xrr6/N1mRLW7jIf9sRD3/
FMRPE2PbMK12oam4uCgGlQH9XqEQfg7cyitS6J++aOgHlIqp0MB1h7P9qRApkZdMQp2Zb5jRVFbP
SufDywvkHBxpYWQrMKFhryBvArF2zbcAuuLbT1Yw+LL9QtQJMOXc5hjukynW+r/EuQntRwR5/fOq
s9mF2pZhX9iTWsIZr7x6dZy5Ck1u6lPG8/wprnoJnx0Q5e2oJzRvwPQKfcDIsvrf3LHaOn5N6YVD
GamnrZtcQhsG4vcp6vpT7HfeBlzuXQ1l6Q/xlexi1943L4PU6S+Bkh7khFFys8GSi9zyCHrwVtDu
9qVw7kmw2Kdzx2PUN31QUEZV0aa03H7dG+wyijXcBZf94rAphP5r4iRRwQqBubMTrizGwzbmvKIS
CN/uyTJMXxbT98ivrss/9GMX9KQ4ejW0IoLeQuTgY0GwxH4M/XXXQq8ExzLnf4e/xARDv+Etzqoj
jMbfXBm5fzUo3vHKzV0CVzkOhG6gSRDSn23BXHt+HcI0iDVRI1ThHe3djVTPL1mQvvHhlWRAN+Ds
9xm/8gLTC04Mg+U90uNhb4kj4SjKELflOEJg5bWFfcVAUWK55PgL8Te90CCTzYOzzZVyZttNpgV6
p8Siz6UHSQLBmAh18v1XVI0y+2SDNVKs03CjRa8lzOnYmifUf7U5k+xd7NHPtjDYmj8GxLOJGPkN
eT86GdGsFpCB4KSnirO04nz33Oaox4PtDlh/az3ARTd3MeH5J69MCcQNQtcZlOpX9K2JrI6cH+Tc
QKOmaVRVcvBZSVkubAxoLSC8r6UuhaklrXoupSI2CzevGD8Ny+8gdUIKPhE2/aGPk+9mbl9Ljpip
DdIUuFo3NdolPDKpx7hUDnTVyz8ifS9AY5/xqZya3qJL8qaSpNmjqAlciu/RToZYw+txYUhwJN/E
8bQZ2A+l3bPn6EUi57xm4kdk9FvFNry8DVv8GuNTfVih90yW8or2OCcS63GJZUKg7kXlPfpt0XZy
mQWU99HuJDgENX5iVfSLbh2DRosfh4ul20BBEd+diA1G2fpqytEXWFBiZFJrickdWprysYf08RPe
91Yjj+aQT5DkqkIRMc1/NQioLrCIqy1OfK7wYEmgbyBaHDB6Tq69Yy/nnzHVWZ4q3dHDjW/vJ3HF
zEKaMYvkSCbFQ8+fQTJ5NQWcFIHMtbKFUTjsOHZ6HV2/ct4g+byuFwpMU9LPqlwiQGANjA1F+Hi/
W9ppfurDaRJxsdPhdtZiG2jwY9ar3wkEdbdUFX9uwfRx36zpbZzk+MR+/Nf+KLKxgQmHlmyZdoeK
qme1N6Y6d41g3veRvFzj5i8Fgo8pcwtW9UBw4jTFZRNZ1QULVbO695ES8+J+uApAvfUSeR/6abJ9
KouMYWVxZPJjW1ia4tlxtdq8/TcruMTFH4VmeuyTbWJpVKtNyY2EVCTbp5SVFxhOkfPNx97us6Xb
MjtiFbEsHgJivO3yeH3KrByq+JfMTjC9MmBpd5ZOKRV1A4t6bMW/hwuqb/yoWvTQ0oRyTT8QkLe3
9W0skouY/L/AOzA9cO8R/RFX6S4lT1a6LQXv4KF53B7RKG92OL0jU+5Jmkk9t+HhdtpoWJgfhHyt
bSNJVulqPobQAwcAweCP/kYQy0LLRP8yRitYDRNfPIwR/zmJFNU+5cu/ZndFDl74illIpGkfREFb
ButILhdr+Uhgs6N3HYvyyASg9x73XGSKgk/JobCQ4lwTuJrVDU+VGxTAC8IuILBV2qHrafoaQueh
KaZvB3ixEyMuARbeLckCBzp66U8XtGi0yS4UjESj0lKtE2wvgvvuCDsKK7hHccJCm47tLgMpVmmt
AgCkEZQ5uKT6o3W8ogMyd8a2Kcbqz7xi1XwlFbH0ytts97HmD4tdKisPzcBzeByG/vQLr6Dpssk3
hw/5GutbWhG1Cw/6cNUf5shG5uTOZNF0H8IufD000gc87tms2KaKBIDjdDtEd9JEqb0ggOZGG3U/
1myUfSTYsnogEOOEU5oXKZO77J9gtMPogAJE/cGNEMR16PlSqeBEmaLePwkVHQJER2nEUZu4qjMr
hurDmCSnXfXg/G7hmN83U2pZw3SJk25zLuwXW5NXMbZ7S/ZWiHL/t5BUufffRXHd0rHbKhq505ID
QJ6EabWgLmMnyFzqQX95JQy4tAmCWQWyKBpXxclLBHbXwi+ApLzNwCExpXU07lNDARYj4egTgN83
kUprk5KATHssJ4CKvezXoAchM4AfYqIFufJspq4wgjc33Cu40aa7G5h0s1ZmHhEh3yms/Ljv5Asy
DJ1KyAnEsUhJe2OPAfdPT5tl34twxR51VSk9IbKlr/gizw5fK2wGuN5PGtAb6eU5X0k0GlRjExxl
D6otztGncXXFsJYBp/NhUSy9IRcKGPSHAJNcdXHV/rwc37ORt3piHH/AJvXhBDh7NlfnHgKoToi0
I+HGx5ZZ4PcJ4VnYc1mp2NNmyTZfY2YEKD617oCJlM5H/7XncKgT36XjFC2BVN/UWElOpTLRb6uz
4c1uLj0JiR1SL9BFdRT8PFS3aEDCIlREEaNnEuKJZelLRQr9TVq0WfLxsa1NC+R8JZcVtPCE8HVg
jpMSd+gZB58Db8dPmsqDgvc/s65gjSkZL2UHXp2kfBVzjwUPHyCOJgA0tq2xA39goM9X92Ik6jzE
YAc+i3xvCsWJKplfJLvbMQId2E+uDv8MFiw0RUTd/6Cee9EuTGYHo9ngWerT5qavRdu/Z/bBYpnr
StoXJGg19gmYqnxBcacxXcq1NTRp9z+e43+JXFfPRsd8nzIykCibGAn5CgRC27l1MCOfttLNtr8C
KChfI2VbZ97lqFDRnG8K3AnsBi3Ma7MjMHRaIS7wHaX0ebEn6bBwgdjLGgo8abj2QLP8oX5oQgLA
Wa0+JQhDN5XuPQoLbSAPeB0DbGb7exMfYNzFa9p5fzIrag7K4miPYTkauT8C96naSBvWlyPo/EUp
LDfPM5a9uIK7HYgtcAkSoIzhJJbf1ToVmSszTZXYYD9i26cjgQTr8zkEp4cajWxjpaqiSYNi/ML/
EwPeDj1y/ogsya4VAPP53oMAn8CzoejLL64kQQIW2Ug36RzALSNZTSn/34avx2SGbaiUVLumG6TR
+ecLGJeDnApaUXlrCLxtT7jht6FsGP16zHqKFEDgD1DbWQ6MLZS5lUXZvQLmHHmn5MFy/LUHFQEx
t5CdYJuzEBsUAYMq6VJXKQ/VCny/tALIvoDl7nKQaCJkxJD8lLJydQ8OgztnqTHAJwt1zPTqorD0
wdamfSIrQQPpWqpRrnVm1U+FTV6ZxI3zGPGCZrUGNsnYsqagWI4aAjq6Oob2YFpn1yjQgAtm0S2x
FDdUf+lk6LDUBBTCoKgIUkNc7f3yk2d7NbAhynXAJnaaGq9PWN+6bCLTZF0ECePVTFM5E4nK2XNR
kmD8wDCnambzfWg6J8m9F/jgxVNYcYhYc7jc1j9gVlknykHp3PtYIku19gOp59oPeGiuqDCDFx9o
PmA0w1FdIrkip9KS2QKk3KIxr/EjzJdCt3dKSZykkbR2knVEShisDVwnePVzXjpLDYSw3zdHdrsA
NTZ2pzj7pyWNP02mqKOT/91kZJQDpc8leJmPqvoM0IjNjR2WocjmxMNdhJIX355yeJnE5tjdiiJX
eC0f8/1rf/MO0J5spAbbR0WQOdOSLi2s2amjwSF2IT79+F/cI4sNCmX7PGpdo8FB+Kwt7rYy+TvG
KSB8yoRa6xEaZynyw3RusQy6zzGqy+L2LCLTDGXjxc6dX4FipQzD7kov3RV2bva6RlXvdvcJjQ1/
DdQIczkMl8muy5PB/SKRFsF9/L2DcBgLF6nt4BmwQR6491wR3HGxy8W9R9Xsz9b23jHhoKUJGH9H
amUog50KZzcMZJF8NozLQJ05JkS2v1KqdPI6qxr52QR4LZQxNcwUgq+x17aRYdxGo5Cc+sD2hDzM
ox+HT2wwjlJfTXBZ1oWYCYVU8hnzQhzCDqR1u/vYjEQ6CB8uNHx4h4XXYcpBWaB3S9ly6OqsehKt
ote5eZxJ3kE2PWzAsfV2nt1ZOGObZJTQ88mreaOMV6kiksYhhNnFlYZAc8yp9PYM1yXwBT1uaVlS
vVXBVY4uBBNslIrxhE5ProTPZUJcNCZHugN2X9gpjAmbtjKAVV6beC9VWq5aPLVs3Q+di4FAupxf
si65Q0Iooa3gcerfeMkAzbKwqx3TE2y+6MRaxO9trUE0N4bmxu4Z2VkGKHuRVMblBjOgPv5hb3mR
DgqwkEK6ij+xTJYRpmu0UbCwzIm6m2v/MDdoJfDawqtaIEQGjRpz60ScBvss4MB483N9wZtui7UB
ceVK/9V1zTHYakFnW0FDg/8xEXma+HHvilCB706kSRJvbrUlTRxtksIlPcR1rUpfspBp8xjfG0aI
yJI4k3U3rYnskK1GGSS7n94hyEWa5kLkzjxs4jJIGjNSzSFgWZFgyjQcUk3K4itiYk/kaEKecRky
KAR2OWJbS6ouDGPTaTbGhLx9nqVqbJN8TPAmqlDUf3746lyaZs/+l5SyjBIros9QKu0jAfXVv8mM
l6fVghDGosPOgL8C/9HeL8hFDsKf+Aro85GwqE7LDt4hFbRFnOkeVD2SpHnu7FRBBla6Au/9y+PK
wlNINNUVWY7C2goPVTNObnIMLC057FRwvushU4DRNc4f2RTvmNRRIaRPd/EEo9VatFEAp1RdENLq
CAdx5plUk2RB/PHgZIfFTWTbLqDdEMjdkkpEcS/jVBdE7yqrdAu/dmLFWsFNfOIPH0bhv4zJSBIe
P+CQdyAT0g5v0+MWevXCbEYpuZv0kos0XUAsSkyUQUxNacx3fxkhtb/t1di6Rvs49qgzc/7eFT2G
SwXP5qK1mf9dcd1X3yi6UXgF7ry2NScaOL/WxVJxAsgKCLo/L/q9NYK3HOlkSg6WNJBeo7t/rawJ
cBjeLazkE+UhRLGUUZAhaI1oowqt1YoZmzgPICkY/4YtukRch2gIyJKxEQCW3wlnBAQaKNvY9kZz
y7whAMGv8S9tA0OKTSj65CkbyOALtcpKmVnnzpoBxXagO02K9W+EGRXCZxoT+hOJs+VpX+PiMi05
a5MKAvUy8+I4Lolgbi+MOHECv+YXK34kFJyWtohwczMssQghpY2kiuZKyhcXbtVipFkqX6GW9Sz4
Cb3YPEm098cmSe0SI4JiCn6Idnd6gRhClqDNpUaRvvh/zleuA8Y+7laGpWYLz4DBHmcUiXWJOaHs
tlySLJFMn5X1sf4ZlrKHt9jV8Lux2DG/5/Wwq3pKiiLswgRQbY3caShZdYPMNFRlTyUavWb8Cazo
CyefSJuyEWZz7szP19/enDAp9ZAzU4t/0N9KfTRgJd1NBbbPGo6Oa8qsqgGTySNm8T8OtRyrMjj1
zouatcEfp/P226cRIDVBLT4lCMGyoP+CDEEU8VWDQvJkwEWvYji6fjjqilwHmioOFh9c0Kncj3al
zo642anjTFRl/XC90DAh4PMW+0B69dTJLWHNF/KB3cI75tSqdivwypyO3zUbyiFioxzRa/vdIigt
S/8cJs0XQslzr9uk4IB8XAv76sar5kvLkfz6M7u3R6rw3GavpG/Acw1Gi1XWAw84fK9syNhUP0Ov
9EuICbGhV1Kw28H32vQ585fwyMF0LjnAylzhiAHkDY/s2244HaCizmNdn4LROVvOi9ShYieWGEeN
Lxs6rBLaNZEvTzp9/wyLPhETGjn3IWGZULmEoivd2V7bnYSjqFJP2X0t8mGQiAg9TiJlc0VI2RTh
zSCYA8gRHAHfyENONF4vzqkLhLmvH5zYQSVwCbPSQFkd7TUaWXD26x2Zd1ELPZavlqMys2Bss+sx
0rQ+opDY/H2pdC/LphvuRyCmK6kFKnVk77yri0/Y4lbQoLBBIe6SSEjt+lkZtIDt8zGRLucVvpvT
J+VU01k4bgIGn30/fwJDtsdHdmaPb8maAr3QuUrdh/7oEN4NuK+0Ze9mGpYLP+vV5OiDsAH2Dpnu
/WGtNCx6QHqsvOcbWfOvQlLgUG9fGZ1CRYlEXh++NEbOG6C5keq1bfPFuXeRAueSC1PaXufTfQrv
kLcco3JdhkIK1uaTdl1qgIxk3Jf9ddYLvcD6eOlq0JzqLf5c7G+c4lKcQYz8EKc4jKCjgHnlTBkp
q0T/Pw+gPNU9ouUinWjs0eshiMMKjdijJlxVo+PjEsqWxYSDO8tiiWQRM7xDtPRmJ72TuIBPhv8r
lVsNZAGtKfCwC7GgfgkgcgE2wqBfoTqkAPCuNTRwPS1sI2Lsn8FhDfqNUsjCd7qf1MkTi20vLpBB
slYzifOYq+6EJk5+gCLcSJyELvlp9fFpJFMyvZ6L100z6SLkG0b25/udFFmUPm4tINmz/DLATCE5
UXcZjihvw432IXNGyRCSh8GHyn6TWE4BVHL63oTu1FPt0Sv+Ew8kNTUNM93bWetiOflLBRIg9vas
dViIzKKN9zJSo5aehssbueLATbhst2v5kOzrdWpUNN0Ln/uOlFjWKxCYU5Z2WRQyHOueu5N+/b1B
kAsj1wRe3+eIA/0vyBwpYTBBC2N3wpDfQc1xy/tn2XHMuu/u0u+wK2WRP0IYY6R8F5rQiucAZ483
5XiXG53puw55BVDFWUtKCBcz6u4uIf5uGLpZ6JNyc7cEVqTQ9KTIzRi/L4qhr2mzOm8591HV9q6r
1h5c1pVECVLEBRvQ5yDkFY5ZssmDemhAp2xpSw2uQC9+03dQYnb0IRJgDzZfCYss9yEuZTL2+Xb2
8zWNWs+eyIwvwfStoiprzQSuCo+5iQcZdtEdyxLifOUIRTaSHkuABAEiljiz2jYaDTQLdyahyqh1
q0FuvR7fOyu28ZjG6n2ULUaWAzIqK2Aw/B2hQQcEk7G+GCyVoUDjN49vNWZgAMSiUQCbLVDHn5u+
HsEvLB6NGvqCFnxBB1nDhvrJg0aTcTwsU4ab+1uJKBzxKmXTqQNvg777vg7VY4QGA67ZWYCB56IG
IsmRASm1f8AugvyCPP8DcYvjpe/RF5vXrhs55ycevZ2SocGlrNloBvlZamJgel9CqrVaerh/HYnJ
JJCQBduMy1LSMvfyl8AAE9XQsJi6zM9Q38En5KAybVtwc+GWPIyG+Y/pDNZCvwvLfOgXFbWo+kGO
YIT5Lba/xgYfjf/Pns0GsLParQvZJ97J6Tnvfy+LHsM+We2zC7klVt8HxCwjnmSrB9+9y/xhWtQn
tXLjnkdDsPRWJfFUWEsTBXRY4Je7fjXYhXYzu+PxOXFEuYMZxPEncm70Fq5RlsILGUvTroZap+8d
zcFBC5bXtzDT/j0l3bXQpuQUwLwUcwgur9C4RfTdbzQcnk2WH1sNk42YLHur7keQFzXHJV9meh/s
oaS4XbFM2GWSov9djgc9+XrTtQwsOMhhkJ0j1SRJs4UKRxkplCPXiY3+9t15W6fiOTFp9x2TK4Yh
nIL8slkWtqisuu0OuklyykHQRqjJcoZni3RJ3WAa0CN9/ZumnKxBt70Tt1oiXlZGoninbHg8WcGH
ceJlJGZUJzJKaCprIFq4HWIqCiYqvqyexPSyu4jyZN797aCXpWvoYxnf8voYir9fXq+ukH7wboce
utVodklXtw6fkYzjaVZf/HSei0NM4F04LsJEm/1Q6PwAs4od8kqDie2yfQYaNzV9cbpwxuFe6uBg
uOntpUFh5XB2g8eXMeDT8Fn+jCk69Ih9y68zbBPu+qPSG7+FOyfXF+59TUqh/BnaqVCT62e4uJI1
OvHmaHV2I41Ge+c9VogRTBKQ54+/wWlTJj4OMmAJUAff0ZLT4YbhdHD4SKH1cLNGrtDghO2Yfah3
YGVBYXIDPHqWJcJme4KxLfjXY7ZC0n2f3VtjJVeVbJ2oGBXqwWCr3EcXC6kt1YxNEuZOA4pX8Z/Z
SoYC990hX6wP1aAJ3beQfcVxw4GYMlfjk0Qg/ETKdKWcOSM+es8XqDgLyvB8x2qpwtKuWxv1OeN0
Gk4XFnT4KuHYtC0xw3PFcv8+GavKSVSXwnmQZDl5q4JbNPhGkZdIzb9U+z1NuKNWPTmjDrTs4t8/
jtqyIGC193/7MjQJJx1oslfpQP5oLKLFcDG5+bW9hGV0wDbEyD3H0V8j/Tl73eFe5gHcHKPOqCJT
ZfSNMdkXRhaKtpHrZOAxE+FdBvEK1SAl/ETjPxizf3cpR1zl/d2EFfMZzIgwtb1yj7rmfB62PHde
YpYXJcBo3h9ZNEkzGcq07rNz9LqZO4nVv9B0yk04dLxYA+EjUaSL7rLJlpYL5YmxhZXH+bu8bBFS
5isTvILaiVz4twQbPdPaUYISj+2qF3GAGvSHxDFcnEHI9YQXB8J1HDjVhXaCuVpix8VpC/tpBoGv
45djpVTI9R+ujq05bYg/LemGCkm17128fE0cecRqR/uHJizepJ0YxgNl3qnWrAwC1fotHo2YGGSd
ykqcaCTNpYp6VkhBEylD4exYa6VCqMLbFcLcH3O6IRkQzl9psQ5Ycxhb3GTKyUlCZ8G+jHLc4pQa
aH/cjwxP8kZsXBAbxpZr11LLpTloku8nkxHHdY0Du2swKPU5dquSazcB81Wb0yxO0WWmpZCo0vVF
wUE807e8tCqJBVvuGqVQk/JRGjE/vMu/6CeTDu75t8wgJ3R1b9s7BPC24gLq9GLAh1Cmd3e3Py2e
RDGeUynHSeYQOBLjuMhsv0ALCfLrVlej6059Jn+FovqXP6YC27/3Vjju4WuYBo6wANUBO827ddug
VNNUYGeCk7/R0R/WlMKQ+uvp5h679M+g0HjBVqJWYIAqzTfrE/UAfm87UOWEJpp5ZP1S1cScJofD
lzyPYj98ShpZxn/4idVUZuQj0A0YMrb/uIjfxKlzteH9pGIKbyn5zqsl55tO79JasO9wHnOY+x6S
FOAV5aDHFtENCSin1hUANPznpHk2T7E1UA5nD5NBtR5dNu2+EW8ASnOuSNTaarDbghPvGyllD/JY
b3LY8xxUKvBrGpNrrczC2JHLpXABLDrhvghrv5+Sggm9gDd7Q5An6WrAnvE4Jsq0APHk7Hgh/Uae
/mhMe33dLVKkx25fhdli8FFdNb8hneDvYgVC/J4qjtcdjM7hkTLVtf5YcA0D4/r7FcPk7v5hf7VM
30i0MnZwSXBUAoxDL5dShprzhuDLBfFrZiSK8RRO3N+hpjsURVZoAZNSIoXigu3DBuIkjItk+MBs
jRM9P5PJ2EhS4bQaPyfF2bDYkaEQ6JL8dTBQACh2OYLf9VpeuswzH+mFRZn3dXc9UkbePNxiAFqz
LUoo6YG6ClrCLCIkFzOgOTr4VIaMjyO1n5hM54Fq6P0QxwMSs1UUoFybSByC6fE/E12LEsFPsiP1
ojndIz2dOs4cB9IoxcYjoAeQ5/ko7qxgglBwYib4DNvaYHx5lvaj9eQBJ8iB0G/yJWdMDxrOms/r
e+5FatgpbEENj+A1FnTEuG6JCid89OI+8f4hQiNI32kY1jblNtcGQ5Nz26Nu3Zxr4zZVcf7YWvsG
3kdWcMlNh0QRSwSVPoafK4fgBat+wpzrqq0v7ek1Zwycq5Hd5lZ+1SIAZaKTU6aUMcDDI2Y3HmTM
WmoWX99tmkJL7dswPY14xccN8AsV9wcm32MaFBtfRQFKtjjLFI3WiSIgn3Aa3FC1I1wUSMHnevxg
RyPgiwBpr4xrSKgaP1dMGQWy9NQxmpmhV9oL+oWoijYJ9kB2CcTQGDIL1RoB1ZuetLCvuoSOFmEN
YflhRXQ2A36KT/ei+I/GWGkfkb+eVzqMCssB52v9Fx6tdw5XNMucHpPb1Efw5wyJ4oIxpEFK7+nL
4HDPmVfM+ePWyN8UFgZliun+/v1hpxx8PGw6puPIVYtWdvukiVBsTzoB/FqfHestPc8I97Vxsou0
6tGuxtLCRb1VdR9WG+zCKVth1xtZVpq+RrKB6MyTW1DPRVxPI0LZnI8D1gBHJF03NIvv2qF1nq6H
hJuY67Or/6s7LwKpkdFp6XNXNafFYfhXSK33lkZR8u3O/TpSfD7OBb+iu7nDRJFivX1I1zlstZAh
8J7/bbEU7xWiD0h45Li1pw7Y3e7mq2XmIDBZBojgNY7EgWHMLHYbvwH1/9Oe4MdjKcIm1NVD0f/I
4KR4EOzGurjmlsrJmX/3/LDreeLXAzWWguawUCFtrst3QoHUu8/D/nHvL5zQ1x+DahK6VPLQWewG
TmQmyYl+heEkADJtV19JkRkKLN8U1flR1pDPirUE6x9CXqxo65CzyxBxM8KruKXneO+DzIu9XtCf
KmolHEokmMCteT76Tnv1MEPe0HOFfD96BPvc+WMp6aB1yn/gktOeE0H7hTUA1TWLfuul5th7Ac9Q
sbym7/1berVT3mFYtvRstI6ES+2BG43qWfJcfASDC3F8CBqaZn7/btUd/ls25/I9NO4Wj8XR3Nru
A/iprLv/YwttZHMcG9YbgikW0GVxDLvXQkdOlAzqyJBnsdtPlEeNe2vZKsp7BV328F0jeGPX7Xs4
CXDghvBTm+YqwmrDzi4ATwvI32tbHB0dTkb8LKfBFEZwkb8ZlvHcBTXbbKaOW1UFeXOy1YRauD8R
gqb1Zh1Q5HBjulrGb2e1haahWLZao5/VLwqKjqhTxmvZz5jQ6XssJb+q8bwf6SWjWVQZ2mqWKOq7
4jPVLypVSIKFo0M7Sw/QHKfx7F9qgto1YvpZfXSUFNTkF9vEKNYJ8QgXY7qG02C1uqDRWk0/XB7m
pXspMY+XKCVYFSTED2/pzvKYZI52MUYqk3D2Sv9ND/5+r8+1Ahh1FlkoAXBPiDFGUqwONe6AruOv
riy5jta5j/UxtcIRRyE7yz0C9ogJrFSVsCuFoWIUW7WrgY+xz9vCRi911A3uunacY7HQut/ucaH6
nxxfuMDa7d/DPKcW3rG+MmozXu4BpKUKyBO2R2wuP79SAi65fv+r9g0uOZv0wLCFshJUAwssVMaH
AAE4+jDSDvBeFiqDI34VAPtPLvuih9iKQhhoKrsRdMPrzlrdraG1ovR6hkYMxPh1YQ7Mq9lDr3ix
smyfJJ/0I4LcPu+uBfteA2tU92t3W3n5M2B1znAyjawpz1Or8CBm944TgI6QNUft5ZnGDMMoBqvs
SLJmkb1eRhLTtNE8rWiHtsmsJcHJPJPmfnFJr0xrzfyJRtYrhtaIMQCn2rOlWp0wJRB7h49JKYim
ZxpEWpQMa7uP5naX/eh6+UHr2WWECey4eujsFlTBVRlOkWUscPB9s78gTPIWtmpJHxgVI/rrNXm6
UBGZ/9XLrCl2M0C57yVEvMdiuiRPV6VlYch0tkPeqaN+BWl2F73SHpg1ooXJGV3l5RT9QHinJtpX
KMYynWIXVNzU1kSKWsAJ4+rXoMk2scUj+7dsW9QwZej0CI7e1yQByu0I7vsXjJtRppBARtgk8cRD
U6dByguOlQlGqgcTxy2SHC79YctUsAL810LvKsYgFJLJq3eNrtje7Sh+euqDimBQ7NaVJa1T6Z7w
gM0MixKn3Yh6GKHxk96/WTb9phN1x3WAF4wwizc8uCLqhXoMcu8S24VfZePHpbU91ydnqp+p2tNE
Uiykti/HRWSXNqSQgMjZi62GoZO1FfzfsujYXLjiOSUph6wrfVhjMfdyHzQUf24gRkNF5ztoLMiP
Ab7+D5+lRI+ftBi1VDaxt1QL5ATrJOjJBZnd5e4zILxuSbuovAYEsJ+vH2LlniCqEZ23ZDetbJez
l1Y1MxNGjZdH1Z7Thc6dhNDC8WPyKzZ8bvMxGNNuPFpWpVjR1J0kkp+3zJ94wOQlk3Z1H96jC41C
RzGYGEB4Kj8+6lgbgPPH9ts+XRxTq0XXlneF3sNdgMsjZVCrEVy2KwE9LrH4XVK+nZAD8XeOlpxP
qJGrUlOMFAH3dE+LG5w3dWEl0Zo60RG8u2wtBj0PhlrM8J+czlgROw5KD0N9PtdE3DQvdmrtDmpg
eRU7djMlh6t8Ndhjfo2gsG1DZmGUSOH4sDGazcYrmQhZZi1zGy5ArioXw0Lcj1VESHRifqn5zHpq
tVTS9CbqxKrNArJNEDkK6R/okLKuB+QXWdz4dJxw5J7HYgc+K+ACK/InCVYfRGtcXYyWtIAsd8Qh
yK5i0cQgeKuXqVivLfyFzD+3A1VZSiklBayt0f7Tyc4p+KKy19NBuKp2fFlKpsD9lk+0n+41uCTu
k3g1PiPobid81T561jVrxHFQiG30vAO2ur+cw9SJwoz1eRWuQf6BG309YUgJ51AOVLM+jfKMZzxz
b9NiKs6ceXqR6jFbH7jXsUBaPZByx7Mrg9sZDUhGmKrR5JCxIekthCUAd6meJlKtwoTcGTAi0+IH
QMzOY1szjrkv/MoAOhddNBiSkcvCky8gWB+ZMwkSjOApcIsltinIdj3IiCC5yulHO2cDds/mJl6w
DHl75tcCnyek5WEUyP9i240uSUrt4YHDDlzYoLB7e3fVApzKCF6qRJ2ORiiyYVKGmaDjXCH4k3rT
wGGRJCeTQc49vKmZzXGGqmNAyk87JoMdhsMDMGOEYwKOhy2lQIgcKET0s0rPcfohkHHWPycEWY7/
gWIXseIzrYJMX2M+mYeuOXy5dRnHP+Iv8oo15KArfNtjaOigvji53/hYBT0YH1xI/Rk++NYpIUNa
2GdFvhy6QZmpD5zjTOexZigsA8BISwK14SOhbxs2afzxW0vXK8/lMRqtYNKRNE0G/zxist9CrWha
J1Ad0+o3Ag4dR2L8vOa7dG4aXzK/V87zt4qhdlbom/hhc3ZuTfibthjl4+lPVr0ZsW9p8I2cvhNP
63rPziBGHRAgAHsSsoOcn3JelbyWRWG+bQ/zcStsGHUDQg75Lw0z2eihK8sqpvxbkE4y6T8oUFi3
b3IEKJb93FF/iAxpjfllITf0rNiu9NUZDr/diNvlgAcoQrR46dt9pfOPapXvE0MxGs9y3r9a0POb
93Z4XSaXUICYXaey7BgeXd5FCci+56P0CRaELSO3M9E7khtpujZUyT1pNNDPZytr9GAwXqwf6nt6
O+8wVLPq+bHiiywG9ivO9OQphFAMofOvMmyMnd4nt0AlQ7GmHwbLzJ6Lk1cE+JF8tzA088QuElb6
Ant0EF3ANSFKGJs8sIMt4bhOr34LErmmtTxIAplv1rwDq7b4LDAhDhV9LNYpUAJ9BrkvSe3n9hVn
o5jFrdN2tDzeuy2Jul+T1lMfIOLfSu7moRhlN9k+ti8xsO+7NnnG3574HY6EC4xajUMB7uj/CmFA
pr4E62MsBspcwkAJYTm2mG8fpHQ+sMEORUFsZh7TfmScJKpKPXzQCy9Ne4r/wvCeEcOMtc5j0qkD
d2m8r8xdGsLEonqg8L8PwvO6jBIjKOOPk2D2z0mt24L6l/6jkoyOgAZ3CWYu2yUG0eiB1/jgen18
lSL0khX3PmgQTcm06Gu7ri2p2QxyK53bTnI0heqBe0vA6fUZ0wX8kf1blEVYzd1+nTUQjCm69dfP
UIIjJ7c6dqdGt/tf2gfsytLpTzyUdHzVS6Xa3fhwz0kYfY3QoO0TdsnqBXaZBBiba2aVnXWbbZ5o
YY0JP2N9gC2dDcuGpzLG5k3Gu1GPdjnorcRI+R8bCR6xdW2AKpIGvo/qZGyeTlkW+1CwxTqkekYg
uVTqxF2rAlzPQPK0w0EZHcy3KTlT1JQ8LYXNxksg32FDopqHtm3nO3Kfovuvn28NekhIkZgGUWJc
o95LPW9zyMJqdiUJKEq14SuefCyX1B1ftUF4Xu+Iv0XmwyPIFGd+vWbGH6VHMna2uzLSp9bwQ4lI
FbqBvwvMLocnLrae/yEyEBZl2MJQuH2Qk/w/xe24MYFSpxZukEeTEAOPOuZcLurzcVnuHhECG+rd
odageCF+QmaHeDze/bOdMev+M8YSvdCUOHAYzW3rf9z5f+delUIbPNCDqLR7qOOxweJyUZa9t1Le
BhjzGdaEuieY1LfcN7NVRKp8AjA31w7suzktgBrKkbVYFQD63/i4p3w2W0MBv0T97ByJHdeT6xLM
BBqLzAO9ShD7nDEvdI8QC3D7Q1GnnLgoiCsjGuAMvtUUlQ7VKTBPb+LfbR0fHCFZAbCn0wcUWlwq
GgAcqrKC4dQAEJtl6md2+EgP4rDAkl4PqmE8DE4z54LfUVpJ+1MMUQ3hQ/UV3YaBJmEr/cjQ/0yx
tLMdHbWO8JNG52huIqlUo5T4vmX8RMTQLdmuCR7dv5EvaZ0ULbNdV+bna6n/pMsIoBWHcrshmvPp
b0VLzgUl+tpM6iHHtZ2EX3ZmzW0AgveNzox+k3SOu7eh9kTzgWLUBIbaWD3srJy9en3hIam/AowR
we38IB77D8UGPzjBacm2ZG+d1jjaxdFAoq6tP+cPgZZ8WfNO/oW1iAUYFUxRq+zFDMe4ScCZxzgv
08iI6qWuEFpJWhzA1Xio+vkLFvqP1RpAGrXwoLi+tJF0QDE9IAqiswqdm0v4fcKmi3ha/19oT4+2
fjli2DboIBVaZhhhip7eHbIhCczBwj8aTdfmnrIuLyiGvqo6HovGtrTOvih/GCblxA7tvz6tuaNI
xg8cVMzQhEHQLfbuC/kGfbyImGhoFcUQPxc063e65/pVLjinE+HTW94t8VLZJ2/NzdB8eSc2Cay5
wR5S4DkUhwe5XHsy1EikNgpzqK6aGDQTzqLH46v5YXZwm/y91vgyYsDqXgf6Y/baD2uELVEAdfUL
ni00JGi6v0AnKZfsphnwd5pUxCoznq4AsqHUVNSwbJhFPVu6NYbMNPJQdGSiSRQW+20Wk0M8I/dz
ShgKF7/VrkCDvHv9pGywiML9ZtPYZTatz2aQ+gVm+zvrFq/zOp4dp9/lbeJV3w6fnw6gmToZZk6q
1zI1LLQmnegHVqE6LWT/FSchxdmKGhdTX+FVqWvfe1uSlT2hksUszFj2INix14htOkWoR/lgXfLj
OPx+GjOJGDSaS/edQkSsOKAroMQsG1lgfpGWDoQ9q04jF2v8M2CCchXdwUGU+62AuvOeNHkI2gt6
UmFYYKPD+UBtWW8ZBkIiMiWtZV37AuLqEIsDEwjjGvRj0DE6/fknuOsE/dveajq1Qy/+kOzvN19F
Dt8KOqj2feupL/HdlTKxouIcJuQxDLLUAu2D9lOdikIObCOAqewWOKRplDRgjerzTwg7dKIX3QvS
QNoplZA2eiVU3YaSW3W9zaPdI2YCnAdi3yRm5AR0/4idoueHqLQHW9Mr51dcIOHGYGMq++15mw0C
HwbdCWbOZG4ASFZ/jtgSfQD9OFtcRiVk6mtlUxaYYwREMTHwScH/U/pqGDMCljLavZPyJUT1ktK8
g3T7aAezWxf4g6dE7ox/mZmb9lOMbDuc5zVpchd2/v2K2fVFQ7YsK7JyM0X9oxjxGs7Xp/8aGwUl
mlmn0NvjOGWR00pyIigO6wVOoDFC94xwBdPMEZ5Z5h/ucFvYAvzPMHjYV4I9DfcwPZAapOk2BrM/
RORtfCKd9xV3NGJJHbmW78meovhWuwdxZgoOBoIL8IYTc5TtCTEZUVKHNT/60y3s3+eJY/x88+Nd
w3lAPVbRk3RX+cwuUrrxZXoA8xSlqkgvjDSJwaKwX4OFz/9hKxNMtFLlIQlnpwv3aDBey4xvVWv7
AFJmWiQ8l7kAa4HpAiaCiaFEJprMA3LJghfVa+2cajFfxzNAfHCoxBXRJd4rnM48Jlk3uXCpb3ED
nMwsqw0OvM/doFjVmAAn9bDksy3RZZ9c+kJ3pImPY4Moqgto/xVVHolN5Xvi3kZKavGoXpmarpSN
LPbmcEnHKCtT9Zvaiw8E91+tcRiqoQ4WJdmyirxDQb7ub8ryiePdbEGQ/Eos5ySCvth0kD5amLh1
2tuyacdpn6ZptiLBD6eSwBsL6/zZ4BLQlTSPB6qNjEkVwBwtdVcYAkrMr+nEQEI0kOLNk7tRsw6Y
LGCOb0x8kx2K10FlLQECadfHqXth7WQ9eDjDW1UwhXTa4sIoCBDMjWVl78QBOKweLnitBihuBA8a
s3VW5Tbn+Gkm2U/ejhNV4kXVEhfSdkhaUwqzf+cqmOuyZ6ET+AMr9OTdtnu0XApkc86mE2l2BJ7p
rt3QbQK1ELBYvd2FV/Q6ffArCq5eBYdcbtkuVgisomtbPxhKChKESXQoQyVsR2t3dYTo8rOz4l0Q
ZSapk1yrC7VkFYhuWWu6B9FJVfA1vOlq+KYYQx/6PW8AtsebXASBawwVzDKeT1rtDxHHodefBC1Z
JchorQbQnLsOJAuK/aKAXjM25x33DSDKB/EKbs9uv4/+iEIyp0MoRYAs0nOrSEJy4ferl84Iuc+V
di/xnA3Yw/bvGTH2GoBk0xS6Fk7YSW65prCZJM9ghHtWqYZHiTM1C47zOP2ekYJ4KDBD5tGDTu97
1P/DSaf5m5GizjUiUZX2bwKYj//au0TXgVrD4yrvGXHOMsQlEgJ7ZkrraLU8eJVW5u0yUxQ9/kfO
Gbh39KCGkhJc4YCz7znTLefpnA+WtZOfaF+vvLkpq9tGo5H/wEFs1PLuvej7NOmXmAAy+uZ+APc/
GevspzAE4d0wmJq3RSEjA/Yozsn1Ltz3R0WxETax2MD8KwievVNr/jpA7U3tYq2du73//AKn+KGh
P5hlXRn1OtDwhVcx7poTPGL9qtQrcjDNAEGFs4Hxr882exgLSz3DZ+fGTMFPWRmB7LNrlnrv3kHH
kzbBPfMxhm6GhxKf5QB/zxZq7mRnIwtEG/OtnAx01FOy8KfkntExohZfPi9FRzAKvrgboGn/bmPF
6wGBP9yD/thAyVFkzS7r2VludCCykRKD5mO12Wia1xaw1w5TpjAhUGTDjWWOCp28Uj064nJdqjRF
MGUUqzzQMuaJOn1DB+Lc9Tne7ZJ7Y3MdxCWco93ewLEZ44KLfn8O94rbqSfMSzXKfrQcAraTbEEi
ROVkb7xDcVEEqeefDk4OChbHGG5wX2nnuJB/ikJMZGT9wfFoWAEOCXfZRHFjqVpHqJX1nadVS6xN
HeEfr5qzBvwmNul4NDgtY5fcZV2yDUyVkocpYzYkA7C2nGE2Wmj/m5/CD/WcnGd4SDOI3hIdNEtH
/sP1ZcgqkjaV8+6z7Q3Y+CgHcdFECbKBcXTH8icXPjWL+6LBnqB/G8LNbmhIoeIzEXdGY7ejmwd6
CQD7oJ68swV8ZW/kfczk+/1Kr5hJ8n8VfsoOsR9ZuCFgURU6tRXNj7QRfKvEs0RCAc/s3DGYmkJw
B08BYtvk4pOlv0KKEQDCzIae2wEvUkF7CHTDw+euamopVS4GKUeomeyb2sMqohb3yusJU69pxqXQ
sWsaYaqNqXUYZGKZ5TuujsAJdbpDGrf4vRc+aEAGBbOxDkOmR11LDLUmwt1PrDPAaJNLPrxVb946
BucZnieT1HuAO8AH4Ty0ckE2QFU/XzRMItzkSpqa5eRGJTFNUuxk4cAkg7i1c51qBw4kK0A4HaqV
r0tkC80IkShaxxNzqmwx9WYuN67XAx+7XPpSB412WQogEdPkyaaY5GIirXyfcobE8mjINLHBVwVu
73LpkdQqfP0IB1RiQM/uO0JBGQL2kFNiW5NtB+3uaBvNb+KHq2jP67TK4UU2jO958IO9IeFyOWPO
w1jTrIygoVTNPusLaBqmrcf5pSseTiTgOxMNYYDH1RaQlPbkaaSJE34luyiq/wcPEOwpISw+ARdk
MczWx5TJLSOa2157TpNmjw4Iu0iMU9jfSMRxi2ap6rdRxnU/glGeOT+Zcl09xZF/kwlOD55prq//
WsoYqugDlIFdhRrR3DwcZS/ssqA0QgPGNiZJNvh6L9gVMVwDX4w8ec2ceDaw2XxshyxdO1ucRS+y
IH/jM353GBJ0oDASX0WW8ObC5G8shL1l8xgYHL6kALdAOxba/Tt+YM0ZF3mn04yKw0ZYJp3dNRC4
FHysEIaD2y3GVKwLxi2/wz7VFeD1xFPLWySKAp6B4xuaO+DXTT77WtUbjTunoMUaBy3MJEDnjSWv
ykTChiTHBelQUjqoHkOPtSoSG/Hjx/vDOuyMoBas8X6mWnPaIW2ULgGt4P8juIKxCKO7eQPj7bfu
VD62wgZaaVJQwWgo8B+CnfFYwEZ1qt9wZ8KhVKZN76A567/Bc/pjeouQr0YzR9TYdyJxDX0SWbPd
RxAJGD+xnT6+C4EMlUD4sr3fjn0ak5jB8VvDVRheJkANDl0P4LiR1S84hSmZzapsOOM1Cy9d5hDj
VkOMCcw8o2++rPFaB4iJ2pBipPdLkpf5GueeIIP2ebtE8OlEXNAVoq2P7kZerBj0wDM2AFrF//us
/kkOn+HboKmtoZMEsDtfG15579Yjke0kk+pv9ZWN5dX/KDVic+oUyPCArdACIEZOlraAmtM7dTvS
DykSIIaZovAACgXzo1bWZ/bvELUeMiD/PBa8ybxyyIhBkU9wv5Tv34bEwH2eUQaLtaQ+53Rd2UKp
r7VXK0+veDA8t9RHMZh8nmUhXaCh3rrLz57DUyO0Q4aqBQmhGy8jxd/yoEx86LQGvtXpCh+/f9CF
4lvztoaC87Riz9MmySs+g1ESWRii2cTJxPyFH/CFiszOdHkCGHHuN8iUpyhha4L7pFGjmwLG20By
YHXi+Qxgeb18+flRDdlomkSdGuOlmyfZBF64W6ve2rKZUvRi7x7eW87VA+XqGD8GXDc0hPSUVf07
/tMH5zc8JNkQKw9V9UhuV4jLFAyO7/D9zU1YV2vy3sNswMpysFiTpOX+hNRmqipWmjGebiEebUkj
i9P1xHhPIj90qv4jkoYm49FvGi7bu9w4moq1li3CYzy506nP98yjzjywuobP+nBSjhqc75yUgLdp
MhFu8WyC4NdMY/ckbXMRSBz51pXgXIgIfuMxrBEDUN64lnb6/D8brIIaVR/RnCcCIgjyQsriBDUM
HvuW9fUxeTCO2t/0J1+boakT0TNuZ0VfiNG+AxYXYl4/ThsSQYpW2GEmEDtWlpdejSG6Zj5fC+8n
WqMd4Jn7o9038cVuSQHT/BWBTHcp1IGnc3wTDW1OzVLAy9121R4V3yo3DoZ8QDVyOX1S7ZaPzSfy
SND4tGFx0RIZfTp0yoJZau6NpNn6e/dQftGkFAfDQd1IYSJFrGcmT1Axh+Co3CEDX7CSoRWaP2G2
piub041QSjkCmkEOYSOdeod5k/MT2CbXoLuiYflTqu+gT+NqfV5z5ZMA3qFfvW7x067jE+4PB0LL
y2P9z8tymtcsdpFhtsUfT0Go3d9Fhjfgm2dwbpMs4UGFaJq8Byvvz44dBpu5SR0sBvsOUtF5XGhI
U5CyF29kkYRft6uUxmFNdATdcTPRIeoQnMzOQvlogZd7EWmCdx/nbr/mNsBCxBfFbdC0Vb+U/sI5
E2PlMmB56LV1KzjBnpXAEkU6Z87zbY/oFulDF469QrcXeaTOEfU6OvWCDsXv+ZAeMM8gQyLay6lh
1KLWdElUxanLFmc60JYE8LIfppBWGiReSNU1n8USqNIB/OcBiyFzlCXrXK8Deumi7hEDoHNHvGfL
ud6ko7EGOgxLuhDRMaXX70SAuih/xQOs4v3FhV60QrnuopMokaxjELsN1iAeH6OdKVIJkfEtbACL
F3XzxdvqcBt2hBexJSx/R8IeiOPSbSivvPAEG4Ebjkv4zE+V+3Al6quKcjjEOjKuSGdNMqRKo5Wa
MWMEbbqnyMHT6jrGS3mowker7F9GCf/3WEyhmSkzfl1gPx5ZjqBFDT42CLrRhUeLIlhNZjSyW61Y
75S2R9vv0kUuvaU5hb55qWrCxJRaC6tOSbkb4ViNId2ifzpdCmhfjy51uCihq7oLkvgF/1Vr8z8R
nRMbykYXsvLkNfrA5DdLfLZ6frrdYmFKGl2+BGCRwovHJlWVsXk+0lBuK+BaAVUrgHkTVA19iOks
DeTxW126a9jOCpyh8iTtmLoGoREaRMg9QQoUK+hv5gNSWMsk/km63F33KUJPHZ8hmhThB4HrMwnm
SQRxIluww6jzx/3fK2snLYJOfPDxEdhnTVhrl0XYwjOPR5G31GkGu80nMfsXEhYKJK9Eu6u0YEiy
SYYZtA7NFcUvrE/bXLjehMvML1EcwUDUqUMbVJACQmXDE26KGt+NZo6xB0DY+b2hk2GXA/nERVwz
zt2gDPSv4Oh7q33bUIQoHSUhivx8I7lehpBI876gfjLpqfmlTN9WP5IBHJhgq+nmrrip11auHyxc
Hasj23KIy9kHAPYBJ6AaToD5QAm6MGy09UtdQrUYL4/6f208eYUkPnxka6r0LX0CH0//XYP8MkZ4
+yRNevuQ+w58gOW28gAm0b6YfTbrn/kgsdwSPPzvKKuNBYVrGfjuiAspTwGRFNxUmsB0YJ5Ceb1c
YTrauNxxRo3UdC1URW1+PIR2R7sISTuBcSxbjfZtmWJW4u9D2lW24zyxE2iDQ8QCjowrTaGsD4eI
5yqXqtm8v2dVpt4bHX22yEQeu0ApgXpDluE7G8QEgqfN99nC+Pw61MYhTu4pMBrPflahPzGKoaAk
Nt85JeqajIu0V/lfdM73gclPyWdBEHUGMx/QmJrLYR+zLqM/Gkl1NKYXuqq4awvh402nDN8erdwJ
fqs8BkZW/3oOrD0aKebAAn2sBUKc0wMepPSDkpUftI1rE0Tdd3KneZlCOAGEnEul2CkDvWrNa6ia
+RjlKjScKKDuoTlVL/zh4p9gNjUp/Rpj3K6zqQA95kJdMYS6rp1b7ieErRDdKf8B5OQyuMlIWF1t
OCCLjMs46aykVOfbwMJpgZh6MvHJVcZ19DBIZer95eayc+N1Hoq9mqpf+sy0BYu1cZLR+9u1SIAt
Gg8lOFPp57JZvk0/Q+MkdBEJa58ho+6LAUtPqK6mjzv7r1Yys0Rry10gd1G0llBkKMeBlhgrY/V8
MePjiubtLniR8OEbPH9JI4iyD3SwwY8bvp4Dq9rjUDaTAnd2tXIr0VdFyn4/Ihqp0PsgysHbLUZ6
5vLYuGyIzCjiYU3fLgDNVCPJJw9/dsZSyjcefZNXkGY0gKGO+4iWW88bH64Bu0PlUWNOzfj/Hj9B
HbaUX0YfZ4rZoGfNNv64HvPt5KymnMtyX7qQAS49vzVtfm8m2vOWWmi4szm1F2vp/bm/ZIOStSzG
H760xPWT84Cg390oQDtkfhAbRrOjwXnhx4gdLaEfuPMi5b3USlx0OY6vSsppupJBit392EESJw7Q
xVyJwTCSTTfbNdXtjQFdNY8oWUfRndbrSGmOk8+XpVLOvvXM8y7goiDw1b8ArYV5rF9Ncu5pJM0o
RZAoJfJDUzybG113+YnCozyNwrMzCYrhDn5PfDq9mj1knglhkB53kBfWOwc5N+Ik5e3lkr9LKWNW
x5zzHu2H11BGAkG2VeYQaFndteYwX7jjTwduGyDMXO0+xchsAc2jszq3XUUvp4x2N+z7KFewQpyq
qGWXNW8B8ePgc3sLBnZOjWQJv0ky8pH2PkIBeWvF5gXy1t5hy8ZM74nkY4Vk3gZIflfB/2owmtEt
PlGj7X6kx6R+y0iZqakawM4Tk2v86dKfGeKtmqcR1YCwF7p5/K+yiVvIXMb3HoQJrLBStCkCJDlf
M3cLnmEv+ZHBIyabPFIxxYZE/mk7WIT/+aOrqzhEceW6I68Y7w2rQ9GCM8zuXYv+0RaXOovMJPSK
o6Z+DRCcsoy8+uk4T5BgyLSVxJBzxxd/cwaAySbStzOwqRWN6xbh2Oe4YYfa5hEROffpBgXTd9kD
8Nvm0XhbU6GTueysRxcYx7GXttNcYWj8xVXPaujq4xoWMJ+ew2r7nHsr+iU2lJzccTEV+IySy6/6
u+MRDaTIdz3KLKBArcXJOCF6ukeYQ8ccupazjvS/F6hPOPD+HtX0ypNgepD4J1ZDyttoUlqyNzH/
hyKkXR1MWVUY4Uh1B6rGNNG3vsef6zmmhUm9vx3I1TM8T3+KGtRVmErBl4C6Mkoo+rVrWXWdQ60W
0J/g9C1qMfeIRQSP7IfbFiQCtTX9Pr7kotUit9/cvXjgLiVjX5jAoUL5ytibkNJ1ZJFh5Jh3G6bN
cy2/2Q6bzoSEXvciEKlJASUjkbteKSy8A2RyUH83w/4/AX72wK3KNFJIiOjfNLZxXVwMxcT377KV
u/oxjwNL0KayBBVU8d/QKwRldLRcD6nl3E9zp6gfz3hpJogAp7M5z7ideOUlUgWqaQqpkcVpX2f3
80Rv/JRLSN/owUAnR2gXoukPdIOTsP4UhXXdvVXSJmCJZd1XClxt32Ae/K3qgTkvXSO26w/p/uye
cnPiefTKHKwAiLyLpRN2KpLsNfbAI6+OpSh026uX5kBNEVVEXkBGPxqXsM7lOjt7hlWnZnGEyvQN
g2LWjifB9LvqFdPWCZJIG3UXbhc34liPQBA/5oFy91Zx3bHjjreA1GaALujCXXZijEH/Xcfb3Q5D
7+MEGBhMqyn4f617jS+HTfo7J9cWbAC0D37xeF5yzZ2rcLxZ0k/aTT+/q7CRwhJ0b0BhtEyY6xlQ
4eohXl9Edv2W8bAfwUQqXsPwA6yoxPJlZr5EJAwHy2U1XsLLnBqezDq6FZMTzv2DhWN9jCJyXIsF
kjPDfXOozb79oSkrjFIHeiUZOY59MFoLFluOGzY4dULAyO/QKNj+My2R6ps23sj00I6daygTTmh4
TVrk1oI5lhLB/bwo/Taa2d1k1RryyyIqViqJB0yCUcO8VYWAXz+/DLoCgKOl/mH21K/nnLpXQnY6
Bj5B3B5x/0Y9aiv4M9ZmENE8nLW2dkm9Du8YM37/nirmu3SAIneuXqj3HCMlc0TW5RxNrhNjarQW
Zc6oSearV05AOBhoP0U8VdL/Hfcx+O73fxm7DA58Qi+E53UMfFBQTrSQzYO7qGqnndD1PglOT4Pa
T2/ihU2eNJ5270CctMme0abqTl5r3Yx8VaPR4rt4f5fnZC1aWOcq22Efo60Lc2UclR1SPF1O4F01
7S7PA4PuPTfxhhbi2ZBcGQqcx8dJ7VB51daUFzZ1F2VQqbtpk0IeOG++eDWGHbV4x/sZaBmf2E0n
7ZA+soWLiR4qhlekRl6WUtXa6Zutt3XbhIagfhI+nBAZX618GOf1jWi5Oe9D75XKdRb0YybSx8bp
32zfI5TUWgpZ5YUAT6J3d6duchZxByZRmmz5tzaZFU6NmMkEvwyLIyyPWAGuHg69GOwejpFXC2GU
l/+gOzGhEqxnsxD0jsq+O7h2kWt85WcfBMD7FgEMi5nP2E86vyI0jueka/64syJP7pt1fNTdL+j/
P5U64lKKdSb4e7vBkVyqN9ETlQ2lhsRjioZgGcnzMK5QNBPLo4DjYzr6pNvmStq19Aztf4iio5aB
yB6YX0wcK1OXXw/3QnDVNhcKzllwHrw+HvWS6bzlFmEDnxgiZ4xcRF5O8zBQWsYCBsyPHeQpW7aE
ai6Res87VEvHGiYeLtytC74VJrajN4c8fB4sNXfBnhehyHHUNze5wGMcMijVxbFoHLGetBEXSJl3
8QDjJwTixHfuaIHJlOPvnwCDg8ew2mLJTMIMIeQgT2DXA/QuTGpY01GGBM0cWV6vNktHK7EolODg
oY8MHEARM+IMRQn2XHFXhMIPv9nvVL1KEoxyOze4X3Pl1kFzGITHozdJNT/ZbZB1hm/cWVqZ68Sd
YnhmFTTaCqp3sliiRyai4KI9RCyoVeK4erSOeh9XwxNK2ZKi6+IKZ4k7tBuaJ5Ox7cZIJYUugavQ
Fz2m+pVEsFQ4OjU5rzN1vBjqQp8DMaprtnwP7Q8H2h1BTGtsvu16cJA3SZOAM2JqaDwJ/nEvlD9d
2W8ncTqFi2wrCzKcVdDbLk7NiKyKxP4jE2Vdu/dso9HZRPprLsz79SXAesHQgUiSEmzmzvxPAgmo
9LJgn/a3Y5BleNveXOusygSR6ioDUSOkovn5SJIwZjD5f0h0ePqUDDdtlbYoyOwN7WLh+TGXI9jx
KkSE8fLqoaQqjgHKMxsJYjraRfaPQ6FwWcGiMmddXZ5L2BUx5n7AxMYJnjzhhAdVQ8ZuQOLwWWnS
HfydVND2NZ3Mds+5d4wfYu6jbzeG4bRR7pnLO4rj6Mm9s9TKK8xLQXnSd7nMgOF2mppnfjoq/Jq1
MpnYjSi58uwgweRGAviORsT9LL0+o1/ikHUAFvFLbpi4zOp6I9oWymvSiMB9HrgCV9mgSnxFhado
geuM9EDFQLW1J+40UxuyfJ0lnloq2UwfuvpuSM0yoBVnpT/9zlieeuHI3XVQaoQa1OV4Sr7bCMcV
CO1s8xGo5j+USXMdVGctbYcouRHBbi/5ANcTi1Vi6PwvBbkbL/4r7srvpb+90z+If/L3FzZRuOQI
KaDAY3oZb9LiRe68HGgmtDRUpvGiCM/5MLIEe1wKksiXBTk/DeaNWKuZet28J2APgKrJiE5IC35Z
6l6xJxrUNJobB0mbjT75qUH3wWmfPlOIQ0nPNm3rIUNLnUhT5XhhoHjAUhyn/URQ8QrYM8S/h4nS
coFNTpK3SKLira7KGzYy/kgVnvQFSFxfE3Icdu9Qv+3y6JLvGI/bisjSw1JIb10Z4qK+S2FhMacH
SoHPtFckFCMNRtBIVJAq6G56/3wy7qCE9V99G/GN24Dy3SeRaJvsfRXGrt2lcq9XiCIHBALAFMyg
KKghpIMOYDvRJyXysIZyxqPGmk6Sj1OfB3rNu/I64UjvbGg/jyMGnbBzi6NL7L1Q974mYpiVaIff
+2cngJw7Bvwd0sg5WpwV6l/TEVlrphTMVfoT879b7mHHMTjf9T4xAKEXU55bzu4Qo/1eHm8oY910
IQwW9rOyPIb7NEUG3bqntgMEjC+gIjoC3Xb1ID3KcCLLUUXHQ7Rb/ABCHSSusidU1CwKhXrYPCVy
Iwl33bgHFsShDLYUVDr++LGQ4shn+lKkwXEPs4LvNUr5vb7swZEcaDAtKCIn1Nb7HN6V5kHXI0io
L0v/P93bTuPi5WPpAySrgLm4wI+qkWdey3NJpjgKNdVGW7W+bs4pJ6mcai2jSnHlbi0e3jZr3P/z
SUYJgsHhwJ2fkvrLitUlGCJwoHzawsLZo1awVYelLQG2nZNZUE6ZUGWzesSA71VTNkTunbB8zjvS
EJmyyke6KJIbhsPfA7B8ubLquAOk2tsdxDK0UkvBBI9/4K+PUHdldpi5m9NFaSfGYjMRMzdEXZyP
xGVXt/kbg5gS+xQoY6+Exc3qAtgAV51feimj/IoOYRkiqLhGu1iwhrjwGtGfAtI5ZQI8ZOCeNeq2
cbsSPkg6xeUqx90J6zEraT86pgQtcH7HA6/csNPDhaRbBs4gi7qjNsDq5+gMQPfwKoBO1lyvKXTn
bxNUBuIrrQ3vHFC963/JK2MJAhEFwCV7qG3+5AWp5f7UVWCip3TB6DICD1NEY8lnT3AB/SLH3T8q
66pl5GxoFOYX4tWOES+0BdAE726xtFLtDwqkYL0v932bxSXqCp8DliQTUsa4aTaaT8j9hgj0jgBY
fcvHU2IqTIsw5pY8RaIrbSYw4kXBxYfbfNWMGpxSZIsm0+EETW3tOB4PLcGVjRrfEop+EK8EK+EP
FMj4cH7LZgm0SfmmPA5TEiNHzZHn0Cz6WaNA3VNO+rA6Crk117hP5k2+KL4Ybq0vmBi4m0tlbyhr
uKbztDv9m/gXd7un2BSzBLswldZqHUjEyO9CqawrEjLceUmKUht0iXGRh/HNaHJ/coWpmo9zm8gU
F/6ZfQwDqvmz36ETqmsk8vx+BwaA98IHUIiMQElVhrXzOsvlYDB8JKQKKHFoVNVnTPx1mBZSYl65
lCfHN9BEVkXVPQuD/VLuSZGyESv4S/cVdIMRppqJPkC9jHQV1oSXQrpfAo7YYyVh5l1R0wMrF0zf
OJ3dLhBI5ZYlsKd6q1fS7JbhIHss8C6m0z9YTcNRp0S1bx8V+MdGjS1TWKzMLFabZc5RApdDECFl
9YnCrXW9veylgVTI27WqaDg/fgpj9hG5hPZlTUftHSkWc49g446zzwMxEiQiS9ZtupSXa0uzNixs
K5NULAeuI8jAiScNu90wwYNXVmR2TW74lYR9yhSfzCw4dkliouP3vXHpDYflSBMg1y978kKf7aXB
53EhIxzC5Nz8pZnVrv5gz0WEILm1lqaltkL1mofGWXFaWRXjCQHBMTCiRWqNq4XFUD2kDMyhlk3o
bUqvP3sr1ckuT01W+H2Xw2GEy/d2jUfWnOQTpcUZCZHYnkcbRlOhNg6R/mbCWobbjIpIEHU3qTt5
m74kytufPSrP6p+PgRjSnYwMgcKy6V/JtWWmNrx8teK/DkD8SpPktwxZuG+5bFsf8OPtgvHOW0Ik
+uMEpuLx9olFQnjXgib0MTvXmC1W4iIBCReAPrgACdiuWwkyHFT91aWhBVLQtTw3L0bP383tEi7Q
DbFOMc7lpNxxkfXXZ4Itj31asLh8fPGL9DWI5NZ2XxfRLEXIkvwIN0hNrGmz/CHO6wv/kv+ryVDV
puwHAtBfm9LB+khNJgv9Ypd4kK1oFgpbXd6Cs1Agl30e0q23LbyOqgSNwmJhVPoeGadKOKXheh9C
SKQe74LaCXufJ5LwhJ2AzMX7b/jUbhKf70uccrx+EAqz7L8kCwm8OW7j4I06FfaWdIjPuPW+EZTb
E6dQZdLVvsbdPCAzJwUXaJM2eWlAZ7GBF8bM0bv4dCYxB5UMWxAIfe6qoKJvHspMU1s07nW0fBM8
85pEhvJzMp/6rXPMm8XyG99iVi2h+jGxVeykfbQM/pWKkCj9wzj7LTUuU2mKub8cQG3+hZLqNqfv
KWb/2YuYV8GzOjUaa+ZMQIDZ8cDRzfah8Ot3VwZ9ymT+yTiWcgguVAR7Ny6ZNsqNKk9vZcSlnZrp
OchfS8YvcvMixZo66pzZlBxPnLWlMMohdIfKP/FXlB2N2cEKX5ZWJbp2vzPZvz9N5IWTtV9J1ebE
UIJtJS+5JB9fKsyEZnRZQE508o14XRxeXf8frDAzS0Y2+KRYT2akJ9YfnVbcvrMuuf2pqhSdlP44
VHnqDkakeYOcIsB/r0ov8LNpFg+4VTCWsA4HG9zcMOyxFU1MVsv04V5aSGEd4pSk+TL4C9aj6Ovk
hwH6Iyq3/PGQXHgKAQOL2xgfkbZnUBR7/jMAXQEX+lPNvIUiQ41rVF6z3wReQAYyJ5S1tgRvgO0/
vpyE5P3GnG6XkGPkAJrpFzn/PxPKw/Awo+iFnedDh3M15WBGp4+W+IuxZiFyJl1yjph8R2uvBkvc
PfAhoXiYa13xLjJkfQsqZ/5baWL0o1FtpZ2axBNF4HXolgMPdhMOSgDGRBkU10cRYaRp3k9HFpWB
wj8yQyqgW264v8623vZp3pJ9jRa/3z6GeiXG1VkFd20RLSqhgltg24iZqijcaznmr2oWjDHvy85z
funuLXSyFfAkbpFuawM5zd3WxirzyE4uCYOiPL8OkOf1dWcmC774FQfcyhSINX+/luUiMpCh+C/u
4wS9zqlIHV/uqqxDgwjR8Nr+GTq3NFasU5wO4z4dYsW0OPRYazTQHejONSHrZXmnczitBZz96RKw
I980TbnVRe+rXXYyW2wdMLVbKe8924y8qHnfRGi/Yqf2yajz0Rgk6BrY+V6d/RmeHfu8NNnXZao4
hniVaOYkiTPNMRaCCOEUBcfHpuz33U2Ax1X2IMssgdoX/1L5mrFbJtNNXt9jXi68TTw5ANxKn8yn
muJoT5v94KiQc8M3xXcwMhQDF/w3ntL3OFqXJuTI7g4UMZrZtOfByUc2tI2prpxpXupOkeuS8vJM
iHcvgvVf7t3BKKtJ5x16TlM5YNbRrxrJ60YdA7R4eFlSXKPK3Btvk1JGTVDxPv/5cmkoCkLsMYOc
VXlliqJHEeO7b0RQDAzidZlRuFikTFSvAvan+HRz8f06vfp0mxAtCRTtZjVRXk24MbbO04aofwT/
RpZU3ittdFjxB+2OknWyApxdE273OGXvbT4jAKtJb48eBhO2Gj7dWwTk52qlV6Bkk/KsNdxKtujW
hK7wJtrzUGhPklaXiLyAmo6hhYVa83Rju4DKIgenPVLMUH9D+8rnAUtT8WD/gdN+x7UyI5r2syNi
qCpiQMs+QUU1hXg6HwPEUpvaQ6HvSz1e/IpilLvxYQKuLuoMb8tYcKnEJxMYHqmCPmVvc0jxMs4s
6EyxXXIDghYTZc46GJyQiAMHYgZtIfOX+jpTl4uupydKGiEJsUlZNF/GCuYhCGPKoS6H7IIt6Acb
MuTd4CEfeXYqtzsBwprEL2gMWmb3svxX04q5UuXEfr3C94iMU6iINoTYYKsvFDZgAh8uY/umbtjJ
pxEZVs0/2r+GLYE1h30amsuSuhYMStNnlEJhMa+oa2N6b0dqBw/pElR4xYB1HV9YJFehHOZNnr9a
Gwv4UW3ZMlgtstFmfOxA84N2mIvsNkHlvUOexzvGXkJq05YC5tzxWRRn2bLGZbNQULgKuCv/VnAS
fT2WuiQt+tUnXPJ+4pnUUsH5ltf8cspgtvyuCcslu5x6EEYicDzJFgevM6hz5Ao7xcGNvIjL0skW
ksONar4GfOGjEY0S5Js7ziWGCv5BKoITwuAnj5k5D0rC61M0bhQ17DPwgg9bWT+TU/NADA+Jg3qF
MvziTnruePlnfvaMACtr8ZlWZtrzSw7lppQV7V8oOJHqAloxwNe42B3hRjrD9a/N8e4irKB8a1HT
xa+MpztvflMPx46T7Tey8UYaQec8SDt0nevUSXHFHruiCUytAAO3SKJiyVSzoBWrU3gSOjuy01og
PFiyY8sxMwCmlsiSo28UVw0m3D9awAhRc1CxKUKk0v9Mv+WZBWwVwuic2Juoadg5VXzOWuIn4x8O
vx5hyEWWm+QU9upjQAd0/aTtENjCEA7Sp+cvYZ2uS4+C1YD0pZvCU82TKOknw1jFKHydAdEocA7a
bUDT/p7wZiI2v+enLJozu8pqItThMPv/UW6x5FafTwL70i5FIBJRANTh8/7gf31bOSwiivtj3kOe
qlRyu2e2jpbDdE83vTqNlAKRiDqCW1wl8KA9G+kjjcSoPOliIaCvISN91hAKNil2lCuRRYITvMmx
FDKiQ9AqlN63N5m5YaEt+L25sEgLHQzdURbYd62Yv21Ulh30m5Kil94GajlHM6qGHzB9ZYbEweQb
mK/wxJHMKnBmZZBzvebEt5zVwFzHZLG0yAgj2UFTyhbzTdhvMAq+D8fCta+pmcCr3+5KE39ccM7+
x5A/FjwI0V02e1SkcD2fIX/2u+BIGKqQSoZscoTwJ7XyHBzL9kODxFlL+DWW0iNbnvM7pSfpWD1T
zIYnzmOA6ukmJIc+ZPjr3pZqtJGe/BpbNkUCBiD45cgWUClcfaC1CDHogL5zZvt1BTF93yL+40dp
8eMcLRQTa5I/OMfxiNwG0lFEHf1+QyyrMc1cWOv7Mh+YAEy2iH67l3Omespjo7PXhbr/p3SOFIfy
kwU/eWbIwqHn0G4EcdWjWokhBiQ43HnQmEMKHvOS0gOoso+aT9ICbqHD21FZJYejbpPmSgNtwxlg
5UXGhXbc0ZxU6CHCHGp1fPA8ZLJsW4h80JzU6JyTcYrtbjWZPxSMIObRkYZqewF5BYZUI4iHXTGq
LvuVxYx2QWptvYka/AjvH+nv7dP9hq5GE/nOmVCAw4kQneUvgLU8fxrzi7A5SzM17hOhTlTvB43h
Ioss4wxJlc4IAeA2QsZm9WAv1qPYFfqQqwdwopBGIgCHOzV8RjfFu0vbxUNxA+F7HIVjMxCYty4w
TLNQiPTHvHtV/NkgQSu3yvaOVd9F7dz7+rZx66onA21DkschcdE0QJMUXGa6szF9YUQaGCjorXSL
gzSyawWJWkLu6rj9aM5GIsiw4A6hQgeKil8tpTm5ljELEewZCnTwV4agF6OAr35RpuLjvKoEpFQT
VFBbPZKYlicHRw/CLi6ckvl6PHQ/YvU/Mu3NBH5TtRNAUV8lSjJreOXRSb/hZoCZZHoBQjLjmxWa
XvTWIRNwvn43EpPlZqv8jKUm+foddPWw4hLCKjBX3FxEu0tmQkiOKKPUaRf8FxBvoiwJIp/UyMP9
fJCXpsGBPFu42h55cihlezegENGdDnIwF+gWq1yUqyXyjOzoKiEHutYg6bgrPtZvDk+Lj70Xovew
++M/NvKHogtr2csrY9ukhD4uDoi4SqVouBFTrT/K/phto7KzjavAXve6RtWaP1yBqLnzsx8x8M0l
UnBSm5EPOUA9fKLm4XUrINVIyuwVBtu/4yWc0il819oJO9LCU3P1xwnAM3vV7fMZwYRRsy1bj8iA
JAJDXGYQd4qQz6E7p95aazUR0SitGKeiQU94XywED3/IC4QIF78jYONXt+UNfGuEBWpu6xf2gTt6
TyXMUaf7FXmF/2khY99dbzvOlvT/2R8TAavJrg/C4lYjbkPDsGBMp1EbJwxgSIguHKYbFaqJHCNL
TDU4Rn6cMwZhx0R8RHBPptwQWeE7OEfYZsui/nlJ6PlvzuWlheWxBwfRt2r6ptr9CFFmql0AjWff
NTAa4THvTluSJNI1ynZZ3h/uOPSAendwioFkvEYFYouuog5sOldzNWCJH1ge1aYc/LYZgogueDGn
hWq69AdiJMHP10QAgp3XYAhiKrxofnixyLvb9m//8GlMvEPquMnC3wLeYzXTMuBBp1D9inPHBkHu
tKkN2QiyZIaisvf740f1xSKgg0YAwwspsP15UxzxxUbS3z88IU053jEG8JYUlQYOBwPmXM8GzZPM
LKyIg7/Xq99HmWZ2ukrXsPDtcNUg575QvQfmgb9VvDrte89dtK70icTUARnOwL1b2eXZEUVBj5yx
kS/nZEXcFwUmtMPw07183xXXBqz/PJZae+3ks3kvTN4bPaMqtprmBZLeiOM7x2mNq944IW19tJXE
9L28yz5EfsRsfzidb79enURPVwUgOqj5Fu94R2M9XWUyxHtQJsspu+PdeoAYd2N4r6VuI+1uCi/c
2964wQgTyS+UUlDOa4yuAhiAIjfY4JDp9MQlzAfSQnmg98pVc62odHlCJ/NJjWPU4a7SArn97cSP
7++ZCg2p0v3YLnfk9mqyM9r2BQHwlVzpBNrFhuT242Kur+fDZ2mUijoCSN1HkKwYzE1mBC2nYFbU
sejOX3Y1R1nyqsqk/2tmVAlWvPXBz/hG9KhqlGWAa2n6Zx4R/tjxR7xf3ZJfv/O4O8uXesfDdLjq
CeCIehOjnlzA+RtUFwS8lj5TJ7QSKs3HsnnYzAr1qauxF34OOY5dTPP2XSVRAjuP5Oo9i+E+NRed
aYyFHkVvCyHUuctvg/RzJ3dcqGI4qDfjNQ9qY9q08BPPwqE/N6pwYI6T2REih/2InSAWwjE9y92u
YVfQD5Y0TLXIgFYAD8KYS16jAWAgdUkZBj6E9YJJmyf6TJmfJz7LltUC3S8kyagL1grpcq+3/QeV
1jq0uCY3Zfh+ZonZr8tgpvbw8IcsOnxfo0fWtkMsbyePmg5gW2vLJCq8Q7LzkFjWSl/mZUBogU1O
kXk0gxK+YVPTVnNBmUNV64rnWIFcdRGV2ZlAa7xJtjg+aHWIIjomztTK/AtldmztAIhSX91+jzz9
eaKDdmDhSMstzsOpMkUSmIjLtsMMl6/TKKHtd7DnocoWCHS0cPupgq04DbbLSaLhaSNXJtCEyrd1
76ijA+/FiEdtnp4hILDw2GW8PShN/3eu0jNTHxQfpGC1yh0+R3E9y3QsIMQDabH8GEMhPiO1/uHk
PBovPlJAgcKBLW8hV3+vZKW/hfqwClr7Y9EVjPKsXbh8wIVXbGJEnZAT0shkymQav9GNhYO1oGtD
/jY3A1G2Ng8CgA9hexsKWnJMNoSlj/eh/AocBTjmQ/Un63ZUgHxcp34sekQb1h0HOvGMmGQwWBzb
k8JqFezzRg7KHCfdV9Si/iocVwbe/6/GhGj/g7XENftfrGMWy8c+Jn9Bm9ydyy1Js64fpTqHgdrw
p+CNh6ZJYyeyfvoFiJX98ZcB5QV26q6nrSU4Ectyc/TOTr8rC8yL12ladn+NXQYN89kkJf+T9QNh
Qx6Zm4cB0M+efnhFGJIm44BKSIxd68yPFRiPqIlG6YLRE2Ah81P+dz1YMpvE1P/pI/xx+HP5s0yJ
HcAUcDdpPjyU2seQ2+RIgSIpHcywd7hUa9T3xoNML7rZRt6PDO5vM/6UIKIOat4xERkPZ5eIlv3C
foqPprl0SbGBgQ2o92w0nxMzRmuaKsLSue0Hd6OXl8MQXfbEZXsQWXEd22GfXLEj0oxdEmCflYUg
5UQnBPElHJnVtNb39fodnC/IXBhgDncnH/Abw/6bBUZzgCfmG/SnzmkRplJ6nICAXaGxREXdt/8P
eUPjv5Fh7T4vqnECz0781Pukhz6eAX9BdGgbK6asBnLiIGaoicOeQLc+UWrcU0FjbA+tbfVtlZI4
fE2E0PR+ShgY2c8V1Ty6FIZtNMYGanSQMIZiqczNRsuZh80SgUhdHNkBNR9B4Q0ibFiegmQnDnCY
stgWwKe//tuLdnpEVjx1ftKazlJS3+c49Apm9NUsU3sGCEpuLEnRDu27l52hhwOGsqjqhUhClhzg
Ivou1tIaS+FnE+pqUa89zwOcpSXTAeZwPF/avj8NMDGBtKwnq3dfwZApNpXuz/8KeTQlyMZ+FKYk
sW16hGl4jqioBqi09keAIHhWm6PvTVcxtC1oA81RS5DRZX8OrVFYH2SJuv8mfG4RFKCAdiI3NRZP
0q1pqQdM8qyel2+y69bCKioQR8XrVo2hl7GQkkb2yK7wpO1pazzxTk9EV/htgBPTSN+dE6MYujnA
UfOFPurp0Dv1XtBjGLeAiP3g+d7qOzoxbgdaX3bPVeF705bU1qBgfNGIOfi1GWgBFQ/f7Tdp5tfc
6EYTW/UQ0CBnc2ZbQte0H3WREpZmHyprszearUIuEyrILqwmRh+gDYsGbRJ8iCaYWvMNsSNu6J9i
oQmHZAEaHmEs21IVE4G9n6kaCqbPpRxLU594sDfpDUy7UGU0A8+5vznYSRI+iZnShZm6eKqy4iOS
VN2c+hYrSaw5xu5+MDoGn/PkbNT8j6jIXvABLmTvnK+CzXFcIcq+HXsn2AqrKATo23sVn1rc0/tA
IwytmzXabRDoL22IdvxxJajPinq7R7PHYxEVeNEDF3mj+xjanvGqLk0/AH/yjeF4Kyuffo9Suv3E
iUcb3beR2vumf++HLXq1skcrgsqpCfiwPoSxxVJ3vaBKQO8LymQhlVyFOLFCb62koNkg5ZM0Z1Zm
kd0RBFItb3n9EOngt+wPzEvR8Ak2vpXzK8Ng9uz6B8t85Lr8lIrkqwrYGq53T7EDsjE64zEUDA4c
/It5znc3WS4TOHXMrY2lOCmruPTFqsHG1x4bNAg4MyV6rXF/Q6c130crYl3Y29SFBehf0nIAhbnQ
0pasvho5dw3K3v1oUzNL4DncXWG1Mj6a0BumFDcbCA7GKe0iu1YCm9UoqbqMQX8k3Q4bSerJN/IK
BJEU20V+TvnNmJioVqQzIk4dyapa5sv9z4boZ4xOIaSC40rq23ws4vtFM584ngL/7zpf/8uqKgZJ
lKKjzKLWEtWjLX0WbpbVgGFxaO+elP+x7iMLmU/OJZh2iSnjlUAAVagym3+aWzsT7IVhvn9PoHT4
M8dlSL0o401zWr958kagkBDl9jn6s9LwAxbqqp8vtu4ZsejcVc/eO493stKZ1ou1Eqim5BQYFjAj
N+6B7YuV+9CNlhk4oYnQxTRTgLT+AsrrXGOi/qMN+a1ibD1zGW4IefoCECLbnaL+ue47mMA4Njfg
ERTKDXcw2XwwjBBpDmrfvk2pNk0qLGOpl+Khvu4ivfBrYHqRu9KoqbsZ2wsRI3XBGks2lqOWxnZW
CiMiVyxPVVacPoAghC0I6/ngLboHetyYFHb5yYMA1yhIdxmPpNQG39L3pFlJBfE2FTKz2xfM49S0
8s1+PVVvMxViC9hwxpgLeW0PkIrHgf9r8hsdSs9Klh9BG33Dh0e60i1a2yEpQhPu37KVh+rElpsl
xiR0sO9MgCveopfL9Z2czjqpNPUycXu9R9Q0S6Ue59wm1codnGNYJyUFSBDyerh+uqBIA015gCKg
LlJcojQIRJ9ez1d0CuZ2IKt4Ki9ub5hV9hrCeC9s+fahEaAywtVadsArYFCXsp6CYahiOluotxig
n/aqEpXYiSEdQX1yNM9EIkeY6eyw8yVbZshlFAOIpxVlty39MClnDPKxFjGgZczOhKB+ubUGaMsr
idNpoNhg2F5URogezgLyRLdAJapi7Fl2UZewpPHz7ExA0zqMa4H3mOxaUUhuc/ZN2KwiFfAWkJPi
ml6dpizjJ3etB+I9O2iKXuLAil7r189KLXJMiE27MvIdlg2d5nuEStUFe8eCsGUsgvywW+9jaj87
vRGACFxcs2iGXUHm4iuflDRRw5SuF9lcfIgpMSAFxCOh4va6Dao9gmVwN1ABgMQIJeIDCm0pwEhq
U9Y6SRXnILpznF2Ahumra6fOyReK6uk7G1PTepEs0uLcNzMEGOH7jRVy9t36B0w5C1Y2E2cRcqxm
sXu61q8pI++lchxO4ZsRw2bnNSOgo2T6QF6UhvWAXmrMyxqKNtW3ZxfREUWRya9935ljF3DNQNwG
AVxEGfG3msNECw8I3yhSIY3sHbW/zrBj8EBiXvlpOU7c8Bj0zsemxVpwUzraV4E+EvKmlDedJaaz
R3RuPEol+t9dcoO5eDwRdtp9HYGNV2y/xjHt60gz7k0SOJBACw1T+VEdO49LpvDyOgyiSyIk7eGl
wRYArH4jPmNO/b1qZVfJs/5DEAZ7DjbrauOpwM85R6qALE54LPJC3e5s4bH2KcSUXiZzl07zcW7v
q01ip0ySUEe7muuRaHIQZTa9sCPoC5MtALRfFIQlxmktevx0ta9MBtLuhQhz2rikY1CRzImr0OB4
tuApD0Yp7ILHRbqi48UHWbCsDu5mfwD5YKGO6pZODVl6si+2fhCqm28ZmOdq14htodMOux/Hl9TG
2BpgXtfqUw7hi3UKY8bN233/kfiCiUEpStZnxet2LZlEpwaWneNeDnpivY65ywqbELD4l/V0sEvZ
Ui5azJ9Wz8Ugyn8RCW48xJ68cLxyn0thH2RTf3xaoDtQAHyfEDaWkSNbYbniJtA9aC5QMyUNgiuF
uuR7LZ6GdZKBoANpmD0FOH2ncHT4UAgL0eyZ0AKSKN3xVi+cmXoL3+FTd9PcqbYlWeJRfsKp0mdR
3j6Zp0T10nbVc3d1j6LnmNcgqHQQw82wYGLK6T9Bn4GUx2e9GpJqhKynpbbHunGJwU1b8qj2dngg
CtNza6XvlXNDyAl9uLK3pL7TPKMbMw6YgdivNOkX5Iwj0kvI/TpcS6ZF5QCIrddwZzHu/mR9HG8R
YqQLHNAP9cHnvA9yI6SDskrPdV4DMY20XF64+2zT+6H8T0ouSbHHXVD+jtXqRFoN0bUvOfxdgrLj
HBXzOYxLM6AhWcdg6oR13Tod/IATYlNk8yH4Nu+RBK6KbfZLmSMKXUPQOhFVIwa6tXzNHKj2Cosf
1HKqz0GkX8u+PbWyJ4mmv6eq/DSTP5UF/1HMw/tCHlJ52ePsOo2dRvcoxgZBTltB07hfubzYyTuH
8NUtl7HyJA8ygffMIk5/EsykStqLrSM/LPPzMQR2QxwKzbtxy2xRW4HHBrjviJHTCdrSjbjZt6Wk
dG11YzTnj3ckY/K/v3SPIx5t9x7ocN9/h9SHJlEzchi1v44ClEMQwzJ8JGzSiMpjeUFr+PudACQM
g/OfjdfwLIqLF6J6AkUXfBzYTJ/3eWBLQrDMWAX9XbOJpZ5xN6bWkMdN6f31H649cPd/r5cqOpN6
Rlv1OvCoxqKP84BdyMwtiryzqz/L/DKuc+LEy6jY2CAkOOalu9X5xheM0wWVFonEpqZPVTRTY5Fo
TBKUplD73D0SPJK8dMxJbkRse/2DUda78Y2ql7vp78XbVVrk61AaVnFnk+ZpLwAu3rTMnjq/dwlP
kPBvY5s2vvn0dlXMdub/PBo7ttrT/sjZE6YZD+z4FICTpntKVPo+gd8Fi2RGtOlHvK6tl0XQT6x3
b43y3vOY3JS4BJaYMDAVqFjfy1HF3A3iX0IwCeaq25InYo2PgJrL4jKbBF+bp2o+oyZ25YELizF1
e26onMxQ9eEZBPPbqpSuI9IO7ln0zrMdctOX2wtL37gFT7+oxcY/2h/IcLI4ixNSaRCDViXUnBWA
0J/7HYGEcW8POAIOcYSDuXYHCAaNU5bSnrlQmQTCjDyY0Q1RwaRvLAPuozaMCMyX/Z+i78XyKn6N
rhGLxEd09qt1s9WLKI+hSVGj4iMS9k2aLUxmYEayEz28+jVGpe8v57j1bXLfD9C7FhJGzookrYzV
AZB/kOYtULj1e4/F9OKVU9QYtFNCE3hnhuADdIvvbF5P3ywH1d4+HUPV1em7xqDIJJtxy6U77oXB
TfQXIRE0WlmotwC6kfF/+b1JeqBKCF6PHL48stGLS/PV/eiE5rUbxZaeU02eNnRJm52KITr6j9Mh
vHLt/5Y+tkz4F+TNTgxYSdQA19/5QdLIqxtaKvB3nnvLxOWNuVol96/KCK2nvnxY7YcguihXnWq6
k0GzdDj6myALS+JNS3SV6ktOZrvBQf9cfdfExkvg6GEVa3pShslZrkxMj8fPb1o7kKG/RnPfPSWL
2aZmLOXwiZq4DQDzPL8rs3cm9yXDL10JuuVGXxJaUY8/kM+wnm65gKYV1fN0yfFu2aogBSHyKIFi
n0PdYFWFdx/3IGX/v08gqQdjmM22nyNxdiCzbYhPClIWZmSEMEenNOgo6YhkpgqCaTpbc7z+n3nG
b79pY9wJ3h9MTzXMxZNQaSHJoVGu8dbtxBxnMzkZtfnsapogTeP1pIvDppfBs/QH7wSd/XrPCl47
KjFnuVjKcsZdgAo2UzzLOMy0pqehXNfR5IOljCe6Ql8Ge7AykUiF9oXVjv9pUl7eEgj6zFn5v1JA
L9/1c1d3JrjIfWAGhDum6wxdwsZxidi8JtTpauihidl/zpJmMvEyXPPIIO+dYUkAJpDeHrZ5ajTX
3Z9yf7wJyEPftqp6jDHrVRAJlpE3e0LwAIjC5b3fVJxw+OFJ2Ti8cDsGRMCLrcR5vOJr4Fynlf3f
DpLLgJ5O0+8jvsAW3F7Ijj8gJ8sL9gwgnIL7FggnxuWlU7SPpOEbV2U2Uda1cr9zpAK0hh3dOayg
PtmGtXthPRQuWnsgC8iy3sqaLqIbVkEOCuOwvGF2AjV9j4PSk6p4GAcGIZB2Wz+nuRjQDhPDkLFA
5vcrp0l9Msp+SYplCFx3L6aMT3vx2d4II2q3MGGFEGgl8DJj8LA+Y+DLJX1Na1Kbun2yBKTyN1ub
TQXrSpCYO8c+PPT/M9JNhYZxhbzAy/3e+qym1V+GNUPBVw9adSN6Li/HAarofx/LC06EYLLt/GKh
yoo5uSgmwxQYi3ryFtDluLGI5BQVquBNOrjWfcLrrH9Ps4j+o0zqxnuXGpDB8CtoTZfrrw5hjZhY
ubCh8KoSMve16ZnyMX7b6UFb5Oq3NlQkcLWkg5d2AjSBJ0dpZisDmXG978G1Osat5XLC7tXTFUh9
e07vgBSJM6dg85vshFNIlxHRrwq+7YkP8YzUAldWwcku5iScy31T3jsKbm4tfLcp/d1ZdjV1gcc3
Ugc1TRqg8Ri7FozdI/IyBdfx92WSLidY+viCjqdOnkNxfjMIR0aMR5lHLodfY1YzvgudRKqLdAXl
TVUWv/AB07IO6h8ARffY5iOsoqCWDEJJ2i6XwmSUK6hOCGkw8qry0tjNz6alweF4bJ9oELx0hwO8
bfI8bofQhE0OoOnTfPTmFlqmB7Lgs8YwfDxTrKAOTHHFoWN0loSeGmEPMXaT3y2dphtqG4IencwQ
1kownTsBeo7Uw37WP25FRTJQsKASFk0SvgW7XPAbychp8AWYn40TTC455hRt1vXziZiOQK+4jodH
VwSNatcnLPF0xmGYTjnIlGJA5WxeWrlUbN+mJFkIbgKFT3gnz2Vyuh2KU6WxFrMgbzy9DxhW/30f
rEeslEksSOmCD/WwQsswZ+QEav18InwSFd2/SBpKrmcbUDxMkhVvQUKQHAd52GMunb/0+1/s0odM
31Qc5LdtmUY1o0Ac5Pq/Mgmu376QJMT1QMIEouMBHPV8bU0EeLvLALRsV1yYzy3dHbkGUStx5VO2
ia2ZEV5wDeJscr2kVP+G/f+Q2F6+TUeyGgRla7wjmC0bDGHkqzoAleKJzO3kjaqo7mtJsrXuqjhD
Mq0m+R7eeVUfhkkyc8SoJCnKp+wdF3+U34Rk6rvUwi0QbnWrpPdcXCrMhL2WmiBjYJvGjsOTwxDI
rOo5hQ4XOpqJHLQvPEUSuUmoOC5FWWVWece7+DIgg7EQSCyvT+gOg7iJrCl/cijsg44OdqCIQ5p6
mGFpfi/8nIgYMVW+fadkpUTtBjpfUHZteBErl2ruukrkl+lHmgqsuFNkF1SiNLPIbXE+Ohthm949
JNAogLktmiSbG16bkCm2oFF1Ed276YNG3xCdQ3whH+cutiOcOHMGqVR31waUT28r8Kcwvq1s4NVl
PbEfc+cLSsKzbtmlCkDb8SYyOI73nfwYvl9fGVOa97ot7u/hyrO1aRWD5osqmN/iwqj0/digHU2i
gfFZPiUuYpxtKMnTFTqlBm4a1DmCKvfHatuEh8DboS3I1EiXtQiRrKMnfO+PtQc/Fk22uWDVXYxC
6zuO6lzcQCfU92sGP8Eh2ZgZSmq+pRVkfjFNRj5SKWx6yIIeZnWjJC4aea+TKaCzKBQOiXJW6pAa
WcfMyVzw+R6uLpgPWVX8wVAWhVzmVu5E6MeRbCTK1cApUwzhLFiPCpsi1+ja85CjPDp38xitohbq
4lVyU99dvGcuN+Xs/BAu7Tq2AJfAC2U2iEyv8QVOCiKoYlJhmfc6KdRYCQACuLdZdT0EKDRu4f3s
23Uou6oeS2GsgvaKyCzZpG14XX1gptgOUAAl9C0vkUt69LwFoI9A0kWZhtrsOUiOIZ3+VLV4RJNY
HQggIInMsE895qdXBIHXzM3wpYEm179m8LjxYnUClIEVFzDpwUSl/HgcRnc2hESjOg1kpJUw6nnL
cf3vnG5bQDUu1zWwyOYoKpx5WK/n1Cyog0RY3mHhZ3P+qeoymGAb0gszlBlTa5dyVPUS3KwreWj+
z2TR8i/O0wm6yD7Ar7yyhvIeb3GysNDNthnqjObtuzJlbrph/thzgANNt8ejPQRus9nZGWU86t3a
DZtDinKelvZjJZ+NvuBuUQJId0T8m8JDOkOR3BKXUrKh3nlRc3L7YQDW6PWfjNBGChcTfPhyGHeQ
CaENZwihdrFDEVK8i1/q5sDt1OWGhtaHVwxCVbHIa1vlvrs4KUdfY8DGWUSmIFlo+bEwXvGoqQEF
4cuzIPM7NN+xPEpfoxFbCWcWeikV4mqiExWz+vkYd1HnRPBmgyzok1IqoR3PGsTNV+khmSntKnvi
kbfSYIZht9+dV8A8G8cL2hhAudqnEfIm3/I8E/KkUuzQYk70MG0YAXLWhWZV761vQj27GYFIaGUe
OszGjzFerPE5v8T+iid6Yy/XJq3wD8RjzB4kdkztAVhoBmrOXm79Pz5LRBWW60459CTQAtDIptkh
b79xefT2NZ7c1zD5Sej5EWKh5tivVNv02lDohmQhXmH6NgzgSBY0PNRNrOlXjbOAxZqhmRxnuR7B
7AB2xocsce/gZNNdgXS9u0sffd8I/bW4DFfVEmi4Fi1n7HQxVdzZAIHoFPZ1YaCBqqi8GIc0Jm3L
f/0FeWXSRe4IlMO9fyYL6zoWyCOasqVwVTBPlHv3i+8uoxlA/9WC2Zw054CoepYFRaiW2LUld4sG
A67azoNDHJQQg8wOIjHTF05es88j/2L/Cha9eBJqPT7cRrdblnqM1CTp5sop5IChWEwWydGLnr4c
cNRZfoFHm8E4p1TUH9XqaX4lp3KlYRk4byVcQQmY0dcZSSsQGvisypA11JywvmHnQAls5c59TcV+
gwnVMhPlj9irtcKEQKmT4yGIXTgc6eWLUniljOYqzySxyHTSTPKcSnHNyspY1f5F7oyjoCUxAghB
4ffrVrij1eCByphP7DL6axlADK8v4urr1MKwkG9dWaNdcaf+87ZHOM/Itox1SbgaeOgfL51dWgQM
tTqmBHxL6zRjCA3XdmooELmev81AZkzpigH8PZavqROqZXt/db18NPukMd/iIBiBsXVTENK1sVMg
jWUr/Slplm8ljXE9dGMV83HIpH42HmulYkuHdOW5CR05smJstE/lFF1CNRHz25EeEvcxL7g+pZDG
OSmxMe1lMnzElwR2WtB88zokjn5hijApS/jRuWgT9tekFTn9EkIJ2ECTYP6DUxdRdLIPDnC/RgDZ
UZJz9A8Eft/fquPzqYQgaZQhprWxlaJoTcvgQz8iNsGDINqGoOmjAFxw3STqhBcyTAyqCaPCDI4l
F7dsxcuxLW5YvTdWfAK8XsvyyqYt0oGmTPwTOf0kAb8qAxROz4O6GrmuFzrNG/3rv+O2blUiYGwN
k0x559omRag0jDE1djG/k2LcyNVaGiDv38NX/Jeu8ZJSg61ljOJs2OuOKf16cNiCUNSDFXL/W5R5
HfWs4QuiP3IZcffle6tsS4Ml5XX7KsCrYn6MaauS3rELZCOPZVE/Vm2+ipI+1YmTmuyqWmiHO/Cw
WTgKSl97ynztR9gZC3O4zKyunl3azIpETuwxJmWUvblF2tQMytcX4f4+YV+nsylb9RwejdtLiioU
G70ZdbzkDH/tvUm4EQLXp+auPTUor4Jl1BYj7a+jFDPRZGUzaaF4glweQv2b4gF3JK67yiOFurkI
v7ZJ8Uoo5/0mN54IMWxic9oge9P0S3idbdgBaB19MsEd3vG6kz81agRos0xVi8G2079crKHcAcYK
pOc3usY+Cv2Vo29J3tOZIC31kma1fFtY4NOVeLFt1BO6ZQh1bTt0IrPYP03iELNsgnD+9movd245
3Cq8jFOcA23ZsxvQQZC64wfM1oOQdMltoUQRO4qnBR9s31ywSZdaCumsmDr5bgHA6SNM7dloa2C6
UQ7xU2e4K/pN61Tiqx3bQN5k/BnVbvZpwUBVauriAyNXhf4YQvs1dVMitUxUW3tplg1OcBz2b/Jq
PhrKbrF3KML+3BWzf/G43xoaEtA+n8M4qcjJYGf8Do1A57WNHP3Wz8IBSLtZ3zuP+21qYvzchgLg
XIlLElQntf3KiB/m6nTAK/Yl89E+yWT7d6AkPq86gtgVNrG6wJD/TOz2cTpa+nboTP/9EB333Gil
0aNK9Klc4o4Tnmwi7ic+fyKYOrLBweUkBcPjubcdawhq7aSVzE26KdV4GnO3UdyqcVdTzjn3V6HE
HPQL9BUOAWRz0NduXGDoUP4rhizD/qk46m8LvK7uD9iuCKiue3zvuKSIhx4fa77BaGBegUM6diHT
zI0tJD2b/BbghzSZuX1dNAkMGjbPCKKz4Up0ziuNJwWYEJZ0oKF7BUBYMZWGu6bmbofoir4Y8fyT
x/DJbCtXHIADcyAfEWG5678dX4N3/tuSrmL6kyI/Fu6r6WUzNkuuEMkqbD1zb2X5UvuBgCvMi+Ta
iI+1MIS/2jQhcR6BZTibKu6n0BGmb9zwv9Vv5dW1WBFPnznjH3kFqhtrFfo+V1NrMFo9/4Azkvt2
35OYmdGTFus1vEm+2vdXH//RxnIQMl1Jcc0owxFlbo3QbJg1pAiEWZcxFBuA/Id2C+o5wqfW89zA
mS8JYa5kwC2FOKRPYeXqLnW7ar+wF0cLixwy/tdATVPMOaOpxacjcxm2G8fF3edAygouryaxu6mJ
iMvVamd7TGEv/+bh/xNtVtHWRTgtWk6PlfnVClBD5Kjfh6qpHaoYQaSbHQSh2ZMCBOKaqHx47tgX
U7ASc11KD4jvprAJwIe47k+pXoGAg+mrh0EnrJNugybfzdpjD8YYngBgHSDM3jbTMEG7RlDFnnQK
a5XDfm+TdC/No6P1ysY2B9B2lwJkn/3psP9fi8IlC7z57EFrxQembpzcaZ7bO861hgKaEuzZBA3U
hcP/aILekTY6b+HOOyjORtBOX11TOTT4OOKGnKaaSkQObIiiKFbBR9/WkwszcvmMRkaHVnFR/rWU
WeQpCQxSX8hfIuai6Tf/jiHLtmpLjW2agrOC52JxVsl+QH3wtpc8ZQZBgUZNuV19IcpT4UhbEi7O
NTnpakq3UBLUJU4xBbk5W3js7CFSn3RKP5GkG7CilAxXm9fuPHt6TbzPCpfuvoUT//YpSVUnEsl5
t6eF4/DMQ8dMPMAbTMLD5GLWd2/xqjko49lFzzZgUDC89kb2TDmWzUNyQ3oG8gUYH2ApeZHjMwII
2/GJSLFI1Sl1ep/sMy7/fes6Kl+rjsRBQcjfP7c2mh0i6NSEnC4TYVZOxZhB783Pa9rwXMjG9Fr6
57cKytl0QKSiLyAH9tJHbsAEd4TF8TRyfqWhiGh9UXBghDI3wIvNsvBmyNIOF+CVlk/Z0YnGWaE8
Gc96UV/DymzCQNo2aeKGDOGmCm5NMns3rsgF2Q8TipHWJT/6EfzYfY6nXsq6rdIhYRze4imaKFlO
36ZhId5LFw6J0i9FeOSNSLPZ98NbqdCv/U7iOkkf/p98crcEE6dEPlyj0VsckTj54PLq8JkI381V
XMYd+iGXw1RGsu4Yv2sI+/tXOPSRZbt881PyHrbnNDvUBzhr6l0DZpwvYxKVwA1R89vjblYo/zqU
0PuGuaNRlGzheylECLQ0gpQ/WArpTEKJBCZ2RxSWuAt5lveHA6cYkKUdM9OiNYSvnHzcPzZWLzgQ
tz379YFDAWcvXtDu68zsJPoBmlJO+2xp7YOqiHicHKPXfFQ1pLMR9pza5Z2ysQyfFl0kitHv6ToJ
SgnkZn34uUGigKYfIjJLNQybCqMXQzHPwp/t6ynrKudoubEzvht+Kr1SFX6AerJ/Bdylo9eFiT7c
i3nRHR5tTxA7RNf8rOedHwmhiijajPQaZFOOqHOP4aKnu00MJS/PntH4QqaGPoaFrEzBrt6+ZT9r
EbaXfqaVgWV3RkiIeRnDs+B2V04L5O1QOTQ+VJPMBvDzjMkWWr61S4rhvZ6TkSnvCqpCRfN8HItw
N+/d3UZL0JgVo45JPbc93POvOe7z/EpY0vEbtYRezA7HqsVNXnceBq4oYWk9wWgmss37ARMeIFCW
Xui9UXRfLU5sQn2L9/gSJdOLy1GsuoMyrO/73bVzAhBxAAOp8WKqLXsmp/HV13EFfPXAKXvBXw6r
Lzfu/ZtuuCC3j+0Sj6+aC92a+XF9DyhA9ky5GgPacBnMVL6qLtZo0BC6/V5UUoo9poFPiAFTlcGX
lYHWvDnY1FNT7PF5/rmlpodsjDGPbUFd1/2BQYrdekWKqfv+Hl0E8kqdkfj8UewR65NTE0Hyr5Vq
39EJidzd41RLK5YRvxd1sucaqzJQ0ZCBNxiG2NWL9PoMooDUfJL8Bw/qMsP6IV6ncwZ1LMH5muI3
NjLFEKrLC22aU4tfft3qwdNjkHZWP8RCF7QQ3mikMjlg6K4I5g9ON3q/n6WvgIY7RUGKSDLSd0D7
wvcNizzU71Mm51uZ9hQaNha9+cSvCJoyJMlYqGD+X3Bd5AoPz22o4awkwkMDAIxdisXZ7QYQASCc
RNfht3TLcAtklWhd6t6Ysu0JrWmp+h+dBcWgdR3KTy+m9t6mMfFuR03JYxgQd7rwdKUor0mIkE+Z
Nfv/mr2ryqkDYU/FbYKA8v8JttkzVuvbDTjtmFA+OJBamNz6Diy7CoPqvN8m238AhVcXr5nH+0jK
k/2BTIw9HL1MQ4CWSsn8t+M+crnWbvOMEXA957YeklOuNdh1Be6MG7MmFr/UWV0ROh4By+sTufFP
KC0OXldE8ZGzo4BQ3KFR7erhoK5i6hQdKdxweRMt0qIuGpoqlSReSmEN5h0WcuIbYxs/9xiOyUgO
8V13c1DO5Q3ANUaAyfKi/TyZQV+gGgZ053N9g9YEPqPGO6HZh8FAasCtGGbYHHdsY4wlzN8POUeW
aYmT+aOmvsespGercKgOLZXu6iG/BeSA5xIwEPkIUj243T/AzV117tdNXVdCGRn6EeQrRCo9VmFU
pNPCBSiZr10/mUI+pSsNsRgEqkQWbRAmAnbbUJKYqR/OsjfEMz04W5olk8Nqa6Glkv4/dwmT6S5Y
vpaGcKkAlM585bvtr3ZlmzESrVNJ4OIA9gUmJjB4KwvgEoZGJpEr1RkrVJ5bUOxrPn9bF1D0G9xL
QgV3HgbyoX3d2vimJyX6vZRfOFoa4AHoGZ6DZZ3EMgQ8Vaa7dk4jCKeMBHS01LWeR0HPKFcvoAp7
svemMZySlg53LuYCqX6BsZQPIRc5QKOWxkzCeh/yEbscyrqcfhUTJw7F/NouyqpZdndmX4blOAkK
kbdxtQtUls4Su4QEIiy1dzH69Xj+RUJh+0oC1cGAgsPC4ID9HSI5VbpRTbPAXhHFgD9IIO0XQ+KB
8tmjyI2eykDd4YB+/8NcGd25qIQaJjV6gF/niDQNvz1swFcVH8ia/jWT9/HrVwBH2fdY2TG8lYgi
jU/mwlWaYHcKjmxrITQtuBt8RpwWsubs+v+7hyU1vmV3VMsVcGS6RZYsv9wjXSnLasp0czmOfjYt
lXHTRoKFHfzcQeph251wE6iILOe8xpTjMnG3s2nmhlLPXPukHc2A+7uy3pg9ZpWEgMCxWrStodoW
IiVrtl9Pvb+a2XZv++iGK6HARCY23TQFbAO7OqRlE5byf5vKDp5IUW0gg9I1st2805teeSJAcJZd
BUGgiggt/QyiOHI689O7vg01KazWfCr+8BotPAv8zZOIRYrkhz9KqwUslCyDLuNLfBQejlFA0aKN
onPy3CuC2iVLTItAktXlutJIjqKQNdK1ZWCKwFVnjeJc5YG8F6Np8DFna/lJnAsk9DRNXLuY5plU
XwMh7Bc+r5RTjJ4g5yPY+iFJvryiLB6j/OsthW36+r4RVuTTCgdMtwcmv1ubT0Co77sCo0oNnmXV
FU5THLfnjcCidRmQFLHkZMmlBI5IGGtyHYYK0DHtpTyBoze0ghPlOQ8GSihrHnkgSFVEZ0XkZviR
xqTkh7r8Ja17BZnQUOy9yduM6IsnwCHSCwX4oVJLUZ57kXihVM/mCg855Ex/AnAQPz3h6jxxZY3M
EBU2vo2EDzXrEGY4bKvofRzoWYtWMJPPu4sTBBw6pKtqvCDuGBWbfar0/1GbSR9BVB1dbnirh035
lEWeSUpqHIj8dSAtH2YlngCzBJzlF715K+RSq64hhvHdgAwZwNXzxiQmSiPNxTcn3qRmGr/4q8df
lS/SOQBXGmrh5QVrIkOp+JtkqcSa1hK4YrEgS5GLkKtRJChPscryJ8AY7tfHTN2riC6vOhEC+mAG
FgMXsd3uNuSBhU76rinGcSo+LI51djIP31pt1fdcyI0DUqXUiTS2NErrB/fW42mIfvMYjlN/TBEa
CRfdtqDV9VW6i7cDC78bzIDPm+HZZRwVlB1dSMER8sMJYoVItvGGBGnvGlDZvIOCoDu8d3bNwhNj
NIHtoWdDV5vFwgzt4IMLEbZXRAOEHmRluqjjCveXsQZjokFMIXpIrWqEVD7E7lFZAell/nJO1z/7
NmLdHGAqI1o8qDM/wso8quwWUaH5fWNkUvl9ihquqy3GeD0zGAvNcnvba0nie8/Z8vlaLISZLQvt
+eYUKnGAfzrOcqZHxxf1KhZXa8T+puokoezM7j9p1OLvDyaf8Du1tz4fKVqfL3q5nUhOXXLlO1u1
wbPt7oDe9Wsge7ADMqoaTPvA6JYiFo0nj+uKjVC6LkAucez7r9CzjcDOdibFtrd1ehQgrcBfk9Db
WxWnaiC+EfZGep+mu03u4q4xLeH+fyy11oWfxg8x/cTOFoX9lVo3MiYscz0agKqwm4vyyuHwQA7V
+HqCCY91pRcnREkbXkI9bMZO6fRLRVkZnp2LDY//Cvs23z/sFx7kEGDztRZyOMC1rRpwgjkcVAQA
UoqVDBWddtQiD212xXKK5HZJdM0t7l+Gy/eYzVvEhZjy95fq0ZzU4O8ie9p/rIGc+pZPH4U7H82M
ExGH52bHn5YYtku+puytyJ7lJuGNtBY78EoLInPNambpzY3xWOZNduxcS/hp5nr/mMVPU5m5Fk7W
1MCIlCxx77vtNpnZLPAEHdraEYEEfXoINS+0l9MHA8TAdE+s7TtwNjV8ZB4v4X3O5uV4IhQ9VyeL
KfqklryX1ryEPvS4PBn50j9+EojgBpC0b+k6KrTBbWLJsU2SAViAqkr5nlnErum0k+nHvorMc8hP
6+0ZbdzPxKGRw06fFDisXfLQvrHEfaaKrQ/0+WeYehrtppoetsnPxJIoMVBVqyahBww6dHj4wJU9
mVESYai8vVk4E91x2MjPwPZHczEEVP0fN1XJO89qF5ZN/cdh932Xf+Q1tX3E0u2etAy8XQ7vpiiz
AN2GrYkLoI4LgtBBGJ4A0rPcUF/36il5g4AQkx8ipu02qYfybvPGeACKViipvcoJXhf+7wo7pgEN
8LN6ZYLtoNfbsWkWvarRublXK/3I17f+ZqVuqZhXTFgY4q6f3o/Cp9on1lTEw4R9rolVX/jJRUrF
Lgcy5tx4rcW2Jk+Wz23SHbJrVEYHpZapoIFkI+CCgsxBpy9iuxJom9Zc05oMAOSZM1eq5Qwts0Qr
boWc3gVqUUbHRH3t4S/TQRnp59OzSOgBP7R7TgOdgzbc9MALA0AxzdAigNRq/on6Azt/ZaFrlYQZ
x63hQIKwIdPYKHpTrRak9IhvPRxnnT4gKbGQF/t+0ylNRz2f5MkdOChoqr4+rHn1ipUnXqNAXkLv
/Dcikrb7sXo2OYH1O9XAnc+ZdZOR8rG5YaXtAk3YMpOMR7j9duXwcEqwanEgqMXWdja+hYzHPtua
fZg0Bf7iG/glUgX1md28FBRkO/RzyAJISve608p6GpPHr18QJiSZG9N67HPieahoFNf0b7wBavLC
NqmdOsDRKEjY/5mc2MyBK8KeEt4M8f/kJu7hnvKb7mNzz/gmVfd3cDilRlPbDp9V8DUXC1SVwob2
tTbL8Kq1xm0B6eSDACZxSY96q2ocVBVz9i2x4/XafLlcyGbaIr3f+0yghG0Qf70lY48WOA0oy9v2
Tz4qs752jp37Ku8xeSeFFZWOijJaq1UgC+ROBSwqrZ1RgRj3jz10p739r+NXqwdoCYcPBb5vTfQL
9rtlCZ4a4ZBKEAkpqzhHYKKcAVyFKqz56ztUEwlux/+0Bfp3p4kdbmEjYwR9kQzA28iAJPD6E4BQ
fEz0btWqSp6zvNUfwSA0vGOkJ24Uz/NvYYmgQL3DJf2f908foaqnkUPgMd6SEBPYqGESXUgN1vsG
YZGWTAKuq97jG/80sD0+rz/ntfHFUhZDSwuDP6Lu3uPJ+3maUtlyTyc82U9Zw75KNbDdastPQReX
AX6VL7xq0IKibI5ecqQfoKH1arl3ImvnQqzW9iIst2C2M54Q+Tcnx+wD9JLOsbgez2zqlGMwjqks
GPhbs3sw9xGcwu60AVgIjHQrYct3sYpgAHoc5oojdytdVGsN7Lh03fzdJi9RdvO8J+BiTvZxx9Vb
+RE8bvotUY6ka89gp2bBzCCn1d2h9/Y6bv74r8k5V5cJMGuze2llLPMjlZpUABs6Kw4HgfwAvT45
UIGp2axW1AqCXTUKSU0YMuryomS1Mu9lGESJhFlXk4bg33IPsY1lsUXV/ZJ85Qwpm7MkM+NSYFmq
Br0s8V5/ahKxPKKcYaV/JyNo6SS3coCCPGg2O0clMLM4drITinauexwnXl6w0LE7OBg2uS7fh10n
4brsT+QEHGWlMhaiv9UKoQqO9uQJ019nZKN0U6K0sXXDuaH6IBdBxDSrohKWTH0YYx9hz8Aom99q
AozeInyvwPHe2sgLM9BIvCFVVHEHj260PcF2bNdUNqEMo7w1X0X2fqAqRsrTYwyKoXRynGcRajpJ
VqnTAQg+7xAOVnAq/H7Yz+0JECl7Iv8B2n7dMuEhgqnA9kI8HJg5yoL1hn/fkCTN3fwfFNtSak4p
AuyViDXEoj35qdfBYLOIAxaeDCDTePWNspwEIWvFe+2B60Nxp0mDQZZjioNnvXxNW5/2WGoF+4KD
/3Yz2Pvgup2MRDwysQ7e1JAnJrvCwKMpveZZ5QtC72EP/mGtwDe/Wl5boFQ6UcLuzzi6exjwjOwb
XpYHj9L6w04bgKI78/IWEMNauF1aDmNCx+FBAo8l2wstzY/fR6J/zdVC7nElc6SEJJfIDbiHz2cU
z2Lk3M9rnf3VvrnM/wDewyxOWZUIm7twdtjQYpIDIY3bw02Zo8anZurVeyKESfMxwF4XP+Fv6MYY
p21tnkXoZhDE+aQ1x+//canyXjBcAcKXrmPXLvrHOriwc4LmneGPUdk9OqXaXObAxVB7b4BhA7eW
2H/LGrRnYTUe6w/WTfN3yx+wAfEM+XeUGeir9WuPGlr3pp3PODIybloQwNxq95/zoGDi8Wn0so//
UvwLrfE0r+oCwUYEaRCDxIY0Lf9fEzpJVTaFAnC9F6MX8OoGap4OaLhJNvlKv1mMR5wMUDYOpuIL
fHzUg1RgdZkSohy9WBTJnjqybs9dc0MVjp3Dq85RQPIolu3X+MLuNkxnvbBXWp+kzUT10jcYhFaj
ZAhMklhlt1e6QSBqwWRsgGAAKlexWZ/awuQkMoGFo0J+/rdlScVCi6ThHbfFvW+rdDpkk51970hP
w5JUwAU1IYWbWQx9ywnq8P24FIYNzh0BKz8Z+gxqxPz3MT39OLIpw/z7uudi3639wBu5rZDntzo2
+6OnIU3Ql3SLwjp8CoNk9p7Ca1jErw5luDStgZ4YBI3OnyLN7yRELJOa/JkAxWSViyRrelFVSmHd
6eybdO3AqjOhgXXV+NjQ4uAKEMlFlXgqK2vF9cOcsw/9GpqYUh+6bOZ4VsR4TcoDer4rkvBx3/1Y
T8wBZIU0Hed+pJUwXu//0WP2JjeLJxTsyt+2e+QQ6Dmz0ousE/dZqzDkRh/TboINUYpRjJkgAnSH
2cM/mrC3FEdAC5PRMPa/aBL0I2hOfo/og0fM6N9JLSh0vCvq2PGl7Mmn4b7UKPYE+XKK1fh1QtTz
w+M9Wob+DPr44kUVB3dmEYgjkCWwP7a1fX/Y6+PD36i4z8SvFMwhqPrAc8RIrkYQNgJ1OzzdtcYK
COtLAkCPka7LguDRn77oPlg7XlnIboWtRqWcoaAH2nibueTB2OflX+TVrm27KWXfPEmHIXBxorWZ
M2PtAPtTWfjdtObSJivfc9DaHE5Cjjl5TdNMiISQHuczEXaHMOTcNUsXxuB/neCHNmBAXJWWhnqm
CVjviNlexPpG4ncWprHjnJKJpD7R6PJaHHiEBV2Jd1ziFcbVjeG0jfrOCtR7rqwz78+jDn0WHZBf
P6eEosH4nn3gWsRoPmmy2BHdEaqnZYnej1dRpES06w2wy64LvO0dpsNUQyJw2E6iIcDoSZP2JbKK
dho1olnM/PRFAWV2X701FZBW9WYiWgJiM9QVfxPY7Cq04FNveJ5Pen3SLanUZfXsm5xQ/+ZxOUOU
y2X6A4m4gBmWxmOndDlgLf40+cl71Z3tN509zJ2FnZ6cxseZUNQQrGOpdfe91mTwaUnNyrKx4Y/N
KMPviGLTZ1Oxl3Fj/lMYa1Q/Xo40/C03B2n++QM30RjISlNUr34d3an0L4g3iuJFFBKBPUGy1wK3
7KFGPQbBTLIASwsIzRT4epdyOB7vrjonNaFOBWBmUhakpqLqezOnbKqNDqCdvibiJrYgjP+aHd3Q
y0+7QCbUNZNBiBrYACAa5MfWugauuhQyKkh9MIyKFRy1m/aeelQMQwX1TTHQXwmtvIMgQr1F/A1L
MJUnRdo6tlrq54EjGNwwDBHvoYEBqUcoYY3NFq4YBj/mKFj6f2C1bivIAYgxbTdBUETEy+Z2hkTB
vmeen+reWXWymzWcQ7WRFSIVXJI/DCk2AAezk/tDGPkh0Cqzffnm/fS5dt/qtGry8ROUIKWym0ER
WUo0iqadaVVrCLH/WB0jZTvXCE4g7LAktiNByReM1tDhyxQz2kbiPg38S4iowztQGYiRXGkILhJj
THELTR5YisOGqSyq6mlOdrYwB9/Nz/VBFP9rPn9oXCrB+Y4m8FAzKyt9r59a8334DxMzMzUiE3R/
Z5pp4akL2BYQAl+LeXGeRfz1A9O/KHjHeA+eXTLgsiFpq0WqqjPgRFAwxXP43QtcnMdnvvp5FkH4
Xf4UbzUFPqBVQwwd5BFYfVO6W5rQKW9y8wjRMS8xSWg0v8PUPo7tPDp2ba//EvHrcSUXf2/jHFQC
IYJUBoThanp4FEQB0utadF+NI8zmkkFCEZq+Y/mzQf+Rxfsg4nX5qmUSwXM0i9gbIMRlFG4hp7Bg
HIAdz+Z6a1rTwB6DlMhXmcYct/naGPi46SXl8U9J0g3vx+fwhuxMl/WDCIvlVon+jUXecXque1Va
1L1FcPd8MO5ZYGDENAGeUYSPdjRQ/oWbYrQa02nD6LCGSGQ2adYxT4FQvCvzWObeOJDvPyFsC9Sl
rElBUvffK6o68HgQFDE/A7rDzgWRXaLLOvoDnZbMUaYtEGkAchnWF9GdrwZwHORuLxgZXsOd3Rzz
lEzi8sEpKxOtTq14mZciGgI3zyQTCjEFqhzemWVo1PplN78tTHs4Nm7I7/QWCykoq0kuxXlqxl8N
ElyvviI/6pFzrojsnOk/fmjxA8fS9m7SWGJmxv4Shn1kxkTrCYJjJvXCLVXr2oHLXGP9TkNnOSKy
70pfEhcNlkl6EsAbHzc6veBNWpkXouB/LVwthEeqD8oPgWlaJJL7kfzvu9rJjyGMfnxsUd6I7tAr
ue3GhRv6Tgjy94/fuCHLL/jB6+l3UIo9rSLlwAwC9HtluHUzEB5eRs5/htZ14nJBNz3F0tr4nUTg
KgZTTL7T2UjYYuT1W8SlKiGKqzhZBVervxTcHKsLWw/vA+ed56PXBDMKilklY/nFMc26N985fIj6
dWukD5OXk0vQEELj0cvlwms9XVLzFLxz1Ll3z3ZljBT7xtgdPQTyDN9G+OEU38wRAFHikRjmnNol
VkzoqXx9A6Kbhe4xn3ID5iU1J46t+uopAUoy1y+l7uY+wf/k7UPgv/ihrdoZR/CVwaQY6NgdVfvT
TinUJmm441tIul8227OSS2eT0kkScTMLoUy7SmmP1Z5e6c22AzklWXniB1ndZagfivi0derKb/+j
Pe21qhNMSZi6tv6naDCqCbL49o7epXHd+AhMbqhctjR4wmQOtvSuIdd9zSVaTWLIsgIruAGjOZtW
3kShAQ+isbAUk2+KjCpbbqXfDoImUhHxJt7Usj537/IFQqBh5rMEdXDFcMJd0ds21jBXHm8Spkzp
oDrWkJU4g5hNJoXRPJYfJyzRwSN3LkTgnN5Hclb7gR/rP7Qx4rZ8x4a5ltXQLjNslvihSsvjVzjT
55jr7jhe50hWMVBOcZCKMj9oqXH8RoaVzON0dbHOacdVCBBWo82E6x+FgfbG6LsGWat7/Bm7uqv2
bcmU+f8kb+pGjXCUsn42v5aaLKfcWZ913krgcg7a8GmFwiUwnKD9Ax5fEpH0EshrzgXE0zQ7dng8
ZiczZW4egnwfbMPN0/Tb+uVb5lQJ6MGT70yca0X2unU8W36jNuB0ZQKkXL73F3UQYr+xX7iYmAuV
1umGvHz37pZEFRiiAY187jSVPcIMflLcnEW6AQzae/X7X6blt5s2v0bTRyV1j5iv1QVOm6xymthy
oih+DOeJigysBpSwkcDmDc5ny6HLr2HWEMk7PfTuS63rgFJUbXIZDCZ0pfnbImcvSrVqgaRmF6JQ
igODWCP5b9zLNAiNYYkb8vXcOQK3NkohqKOp71L85YvrhNbH0K6lrs1IYJFx1bhU9tN72+u4vrif
I9hzHg5QbUvCbSobEnm2BamHaDA0uhIaL8ymQYxnVucSMDKkRo8b8r5r9r87LAJ7N8wNKqmgW5jE
/T7SyK8Rqam61fdF3RF69qlWfzNE+lduh4obDYto0JZ23fR7BiexlId0LiU1YighyM0ZGnvF/kYt
PixNfOjBPfhSMR1O36JpdR7bBH4FubTh7Aa3ZkIZpxJli8bevsZJVlretCLHZe1pX2lXdNKvtXUx
Z0/bZv1PVCJmWzCBUVfSwikYCu4I1I0H4fmOHl2WfAhsO69r0QFl9hakiinmchh2CmZ/DuckQWQ+
ejwP9BfEBSSn3uebONu8uqKroNtWck3Yh+JHglcEKoGA1PxUVP7tldkJHlWi/WftoaKifFTuzboc
EiqP1hMhnmS0e/SxRdxuVw/EAQBAUFVbCVUmQx3hLly7YOu1aEjdXy/lO718NnMZ4BTo9WiX1ZX5
3uco4yPLZZTjg8ChKukkizD2T23u+CDz5M7XXjAF3S1Sar325TD2DGelRBEiuVgltN5n82efCr0N
6+mgMGQdD5Gab6XJwkqrMyguG2HyudmMhbtbpu7RA3OixrtREZe9FKLrt/3DBu9L056u2X7VeIoO
WCqx+67qBeXpXR8Zvx/BaIYm5ZlXLzaGFx7gbBL7z1V6ASgCoLaR0BH64RYgdfxPHxiea1HyIOEe
alwvLxW3DW7BVxIkIphKzStPE/M1mUmyK4+fLNdMwQs7WLQZXO+i3yrNKxyNoaaRB+9kCqlUohGK
luG4TSwETqNWDAHn9qe+ogYlJCvcPOofZpdJq6xH/5s17IJxPn0QOELFQVdx7V1OEyLhmd52pjMJ
uMixI7VSDQJy6fC+uYKs0WeG55NiVmaELGEklrAVFwoh3SsTq9+6kLQb2gWElSKvZlUDZVeHGqe1
Hlve9EyaPEj4a+vJi0fp8u0m9sdmYWizNlH1P7Ugj8KTHUYTtJb3F61w7QuvccI2pstpJF2WKmd5
aCuylkNnLuXL3VdBCmIgSrD06WB0C4rwsVlWCQZF6xx+7F+tDYjF2yN+7jmo4179QOe8g2uHH+up
/UV00JoHqjdZBkXv2lRmMeGUnjMQ9/SQvshJOHEWfCSuGRD+Vg91aII+By36kUYu4yyJbpdpWIj8
1F+ZTgwPYEIznnDTfs8qFIr6VBsyrSETi1NNoU2wbrvfq0Yt+ynDQUhrlP98zvkjwuuT4/oODYgy
IaUotMuC2hgu/MZTDhjDP6eaENzhWJgKRwfTKS/8A9VI9lvVF1gBnW1EBpTqn+2TgwINTMQZvToJ
JfjJhFHRywJoq94TLyLBZ5V7982Efsf8XE1nuSS7rzToe8SidUJPPCgNZ3lAfsxbj3UC1VZVep+B
co5Z8TuLGLlpTzmjM3dkkokas9ZG/EmWFs5criSzHOsNs+4/qr2XP9lPn96Vj4z0nYuQcFpA5+IY
K6by5a6gamuU4JXQgwUHiQ6+905grbGjiowW5XWjtK2W+yWP2mGc+6064shkGbJqPmNyC1G+dQp7
FUT7zwDnOu+SzRr++P/QrVG8HzyLJasWPHi2GWzYX/LJxlgQJawmvor+Ahg8giAvuwbd63ki2F7Y
EBEc2IkDOYpvw8X4I6M9P7d6TVJdd8K8G6yLEv0rPCMOzuBNeBB+73tQVaIesVlr8EdZlGzJ4K/h
MILF4vTGc/AsJ1Yx5k22s2cMBiwAvKwJLDGrz1/N0IMRalSoZi8LDj+1aFeGeB8X6QkDGNYZyZjr
vTrN6vtFG5z6R2wQwiKKWXbdcNG4auI18MdXqr8QxzJ3pG7K2Dv8knKgPhV7eSdZ3F7mp1+hAnsd
hKQ3I9Xw+SLv+1fewAfUXZp+cycRx4nYNTFHaTpUxelgwNjbSCKQp6JpW0+c6SlXuCtkX7UA0Asx
13bkayGeKLDgDGB/CBD/XYMlIYfki6fIxy9Cd+08o169tO9wwQVLU8f+R+btIdrtA7s9R7/wijQR
b7ovAWahRM35sKyw1lNR94DPuc2065Y2svd6Agi5aUfoIcmNyDptLWaZmF4yokk//eMid58zpS0s
vUfBynTE+VQD+Cx4B8RgF4Ic1BzQoN5CeCMisDHODGLBKl+WauVfanghzHKgJ0sCMTEWdsi2xS7f
YAjDjFrdm0GrwJx5oKAAkJNhjG9K2iHarg95qPkvmSt0F6go0KI2GpKLwwa89WAzo7go23XhwHJo
AGuPXKXsvknesPqPbU8AoLyZ3Db4bpQ+KxZU9hgWYNNgdU6oQbveMOw/pJLbngZaHWuoQ/BOsBfd
Qru/GI368K3GqIu7a3+QNtKigDe5oVYyiUpd2PHO2WFS0O+DToIvv7qs49ff59alhf1bWuEbrcoA
qC/xr1AZRYy6YvRI3Ci/vsX1qMgGqXyPtrVupoVEfpZpKap92KsRRkSVXJ7jxr3O3Z3YFlB88+AV
hxirdnbgFQoDf8APbHoaEqyqQ6JztF5vLOQRfpW1J1gVRRrZb2WyhIMgSkp6jU62Q1MJpDosoZXp
UepEyp4wb7ZsGfaV/XcrYodKa4p6TYWg2Y4VzpOr2MsIaP6/ihlUpMKGXtE9NR0bJjcT4PxE6BW2
DW2rVEPLG/gJLRJtUkvAZtcckBWEGWDQUobgyhLHqQF5tE/KK9kB3XV2FaugOjzhwrst8D798dwu
C/8+EjPHqVVKDRSDwuQ+NxOc9aUsbhtVG3WOX5pPf1LyJMfUycWhPIGH7mYI5YqjU1kqrS24HDdF
tmju8J9BwzUxyoB/Nt/XGo3lLOzpxd0iH2IbdMDjdwSTwwFPBasq6g2Q2g48LT3mAktuFUPodlMG
f9R1fn7786bezvlWHI0QCoK6cjWBCEuAkwv415Me3u8kdViOYjwO7PTmIC3roEe70xpxAduhUYNt
5sCqSaDkJrY0Tlegw0O2kBMQo8E1du5ez1wI37MKA72btmDtY/HAlKtGL8tazRVQ/eKVInG6d14M
m8sbp/eWGc379ZWax14v8r553KQLgg+/mWs1+BBFe/wk9zVfiztBpCbtqWg0iQxKLD4dWlOkyS3a
0lyWcn3sl993KJZ+fkPL80j0Veif7klJJdNLIpj6fJkFlfSzAyASYcX67TmYh2h09+vpowjSw0y1
WeMWTmfal0RM8019dBzZ0BLtf0vbQbOU9pQhjsS8F32WGRZspWZqtXTa0NzSm1xCcJEfgleH1Obh
9szOZJoes1XPWGFl8Kid3A2uDYJNaNFyG7/78e7bf6mR8g1MOnIa0kjVjQD2/G3YplLHjnoRIK79
5yUIHh20yalwZdHDPrSE299/Nw29P90lVQCUxB9uqPP2wlay3MPe8iLmehJlDCO/Rlp79drU/pyb
NnYm+SjowWd/YW8cdHA75/GhBnZTk8q1lx2J61i7BwYUBfZrLodLvGPRr6zYgbPn+7AtTjiwFaUB
pxsmtvIgc11NlKhcuwlN2hRxBKKDuRLcPMHe4pYKzolbhp6Sjs9y5NeUSI1tMT3lpbCoBgzmsATm
WIJLW1j3sLUVNbm8az9UvKjYlh7GOQnN57FG7ivLo+mbSocjDT5nMsA2nhPGAzf77cONhzqOFa8S
r2GtJmCJKoQs4Xye+U2k2TL8P2cIcrb8EZgcDXbMRHQbJZfqH1Gq2FOnnDOUQu6vSpNyrurEGTgS
yX5UprjJ8VhSvRyaEJ1Wah26+i4KOe8OfBpSK1LoYihP+doFIWPvcRxpcsPNb1l+5O8BYoO9hhfc
vwo+yN4WGGOejvGja+y7YOtCAwrac6n5RH9kH2mci+LCiEkWSIojzGooKzUqeVXruPCZ6pu+ffFC
9NIn8qlnrboPHO2eWMpL5qOUUEKwYxPkwVuDk0jdQVoi0vRHsasHL3iWeI365DlEALwHe2Er9Vsp
ThB+DGXZrvpD6VMi2WwUti3SzRSDjBg1VVBbOgLj0jMLzZUBztLzid1h6+pW0nCZkKCFqMs++/lZ
blP7jIqJXEfeYRIq9eEp0x5nQQMQ6c9B7c74dDQMiTdy+zcBdm2RYBgLaGzRul2nykNdDK0BjNaV
7cgGuU3I6mH67htT2pKvCmgqkdtZn+pUvYc/N04zhVwphU+sDLTIZWuYFaRnZEcPI0t9spNBN5wn
5f/YRQyZOT3HWTrE1YpoBi+1v1wQQx/1sSybcbuq2tmbU6dD4vLFtkGMfl+kJ0UXDsL+GCr+SmQR
EmM83m5RjDreDlLywmxzqRPg9wlo4KIjHUVHFK42WGFPTA0UNkGCS2yIz0qziymFQu22AU+9aAQ9
egcDDyziem0OQxPVrFhBUgbSJkIDem4Me3GIerOYIZ1KRfTbIkg17Qgz/vQBvTE6d5dXoxYCY5pb
dsQftOonB5Yz/KiDt2B+884Y+8RZ5T3+kwDWgQvPBRtKJoXzOxjGnhFYCv6WzgAudhDs0EQXiaJO
+MLdi+QYLddFTCpPQGy6fwILc0WDWyjXhhXvTfsrd5yF6tSJgWRQrCGkL9H7kXz4WSPwKEmkJ7uL
5KZc0GTmp3ztiiqsFIhqWhkZLqKIZLItZFlOSznVy6OwZ83roWatWTWvim1ZtznFw51iWqOneZ/5
r6ie8v+QK+qh8MiD61zwimLEu6DW4QLLrk0enaqHswPcTyGyU+oeezkYtLJeb7BD1vAqGwJyXXI4
+2Cmmq5aXXmSg7LOH96okXVVEwvQ/yFY84nrXFVYtVSYVSGwePl7ofS5/dCEIl+fmgl/Apcy+5yj
LWkHUUXggrn/tnPtjGiJoRtay1VvOticW/dt3X2nJfZ3DkyZTO2PokDdRArdSIWOti/7zrsWmHtc
YpHjUyUjYm87Bo3UQe5CZ4RPhSs96c760lFyUBBmUaiDaBTkqpYFZQMrFuVkK3+kjlRRLClX4HiV
ihyede4sEcY2eCQoaYY0wxCbGvOrspbfBDHy3eJ7GTcLsPfFJyzFESi4YGkX46ByVZfzWvYVDb5B
/u+TtTRyrDCMTFzndDhQPfs4UnJpq/w6W5n3kArHxKTTgjZkQVZptolxxL7SoKkdeUJ6j02wgcPn
F0LsTcFTJDjl0Yu6LJvt/6/r0SxRAuwwmFE39l/UfrXlbIjjYrfAjxnNUkX1ypB9eRvYnrB5WJg1
wKj2sykB4FiC1aYM5Spn5m5Bs4uwvMnRaJNxVOGof/gG+zigMPYnzCDGoTUPAtqhAQwD/go+uRNa
FpzZx8WJSMSxjt3v3ReZ554bq1lm9NkQUcLxndMdKK+aPitEVgfv0KLl0zoXSZYaiQ26EKqyqDSB
uObLKNH5OmUnqJQU4rY/QPPC2RLa1ohFjv6BvAnsU20YdAzxNd2NIp2ItoC408X45zRsJOXKWchr
dHHyxlTXBNffCHHl1bY7wo45EPWAhT2h+sIi2rH7dGWgk+paVSS/UJOv6zJenMX0qFAjaRAuavN1
dWkK1jFmj1MPwOiQXbi//F7KaH1PxbEBXSCKwxuVH1JT6jDxAO8hTR8/cUBiNtFYtYZnHPe/U8JG
ClSS8yssAxaVWDTUkVJ+dtbp1iADwimbKpnUs9dJyFRbo6pp4uDTQy049axzdm7h5zQpPHB/uJwo
uBQb1G0Jjgyj7YyZNTLnJ+n70OoJqyljuv92CNQqJryNJ7aH9ZJaQlEADbIWLixJpSNICCa6ugow
WxswBDTzvldoceGLz2vN5TAMaBd/TltmioTlzkwgnrWjTQLgVxzfRnzlOCr8fyeBT+Jp8xQBtPog
oIWRRFtzjohgOCYbsz8quttaKbyWGcxDETUY//Kpdh62JPTUhCWIqyycNB5ZybLvFRzPOyNG4gvC
axj1JhqHZuYZZ+D/sr37x5T/noiEvbuNXRyYUKt8+PJhCA4WpECerLp/xVFmFFLwaKNpcHEveRho
sOQSzJieUMGHYgwrSvVAJuwBMvx1s4U/eQir74UpsxmG3tcWGAOdVHwRwnxkJUM+vG0tPEB5UPqW
wzvxHqbkEknV2ujMstaTuzsrIbkD9HbD7qg9J4jRegC6P0GmjqxlFoJBKxiqm7HViUbgTPd/XywA
OZNtEgwRRnC3GRlxoyYCZQqtgKoJD5k0Xh3Cxu9L6bE/ZQqQUuITckyH0zH7PZatJlbAetWnymAD
YvHwRBZMkMD2RN4wuwdzQr9/Tr1hMgsO0TZjbjAThp0ppmLzLF/37EPMWWchSuRLN8d0jnjuRZf2
jdHOcHsx50rnBKxC8mWBM1r5K99zRqH8srT47UvboHfNeRM0+WdPSIyYZiGA/UWLnFcrlotVL29Y
SHlbpYCepF1WHUBjFK4w3d2qVrI1bUbDPGMYx3iv/VL5jRVBuRE8oO/doj35UM08nnDjj7exPqZv
jpG2DGwreDPzHQVLLjMQUnOJ58KH0l1d+HmOUz4tFN8qcmvq6xzqToPFFqrn/OsUT1p0XWqeoaMx
e1pxGxf09g9DMumkU0dwnTJE7WXy7P3IroB2IWLbmAfZ/Burht4DDjgWOiarvKp/9th0Po14dX3H
Ay0lDA8dOcYrB4qclDYttthpQoXC3egQ9fLgIEOYGEaAuy5+cWtoeCWHGUWulmOYmh03aq7XZoCL
Z6gW8fzMehv4ul8Ou0gJm8Tn1ME7Aq0erucAPp3alSivWZd7rB6WWC8TbQOabydQhBLYKNMp0NpH
z3x54KyNk36Nsx9Q5X2Iq2EWG30d39SvraF17xrv42ULhHZnI2eAhEcpQN7H/N0yCpwjxzT28tTb
0oTnmGYIugY2CvaE+aIYwPMDJo2+hiz80zG+yB0wPm2zgJV/PQEy2LGaeBML2rIx/8WQcyvtFfhI
WC1qAddTTfp9B41rPg0JeDXmVIQOkJIDCWBYkkZT0G2y57nIx2PKteZz/N+FVhk4RedaU4sD9WoP
Wi1xCkeOoLLLmbCv+GGFUYbLemTWdetBfHxGcLLU9gFSFmtQJsMDOjJNILcEXxDXwCovIRD8rnqv
+4fUFUpzju3qAgnftzryJyk2kc6KnHkjZRGYF79iSFg+9C1X4x4ieU1g+ofPeq+03Wth5F8XknwC
2HkQF4apa0y/y1uD2G3mqpNyG5V5eogIZsbprXe4VsiJhFWYcfT8NP6LC6HhJX73GyKmH6gsNGAe
Q3ifJM3zLPDufPtSH5r30IwBFcIrjUpctLt8onc12PCt7YzRwEUwgu5wFk1lbhVw68DuBXq4lTGs
0hvNGrs12h86doquS46vPtqcpdHU4pZxxC8NunTNeQWeBNkGMHJ73kr5iu5OPWBhZKy8lekXZ/ce
7lgd2njNzYFnGX98VctR1ZkKzIb7upBG89YcuDUcG+XC5f2F6iXrjvj6uGEWOSPwCLyadrZyfIzl
na5KUDVrL/WiR3Pmp+r/XTF5FpVcNBZo7wXblKMcg74V58iixYw6xfMhwHPaKpUkmdv6AUKq+LFK
IsFDr4Mx3PACAc9fTWVj1O//xrmSuTAW+FHH3V4eAmG5LdpZ+MY8VpmgE3FtAKFtuw51DawL8TK5
gp/5w5uaWX4I2CKaq4F3bLLioZ/XERQXkiZjSweYg9HrL7mfBKQYZHz2EnnVlp4BhF/Dtzed/zdL
oHP3Mn56hWgV1kpGD1Y6UvgIEch7O5m9XTGqJ3PVZ5rhbTdJzJwIEfXfU+V/OC10Oo40IUrI/Dr4
anaxIE39vhfndb9iRPwVAaGAckVy49xM4mvwxgjrK9DQ47DfIUJJJ7b0iYJDzmZjug5eG+fSDyNd
hp8P7/AbhPhFHp1uGrw5cNy+i+yr15RkO0/uxGWuAKThf31PrNBrH/MbuyYTha/P5KWhHlQnfSWr
yXxyZn4bmtACRPpDyfrC7Qx6NEDLHTTJSie8UN0GaqV50bKcc2qQhkL7uoMJdabNu5ipAPhTQXNw
64Q3/tA05IkBsQVA5nRdoqusKV9CPuKg5EWZFcWo4y3EBbsQGv1V0Diu7FIMEl64bnM54UIv5O4y
9556zpn1gj5Q31mQN45wATOoVRLezHGSoxO1IigtKpK2ex1js40vtPhRGI16uEgaN009M4TeTrpe
mmtHZmbRaMuebmf1LpWPQQVxbmPMzoJDmT20TPPOupppiVJoLNJsTc3oauoGvGyedYq+2QnEd3h6
dhc4ejehQbjhQHXGXJpqIWQNILdG9rKV9X4mdEw2GbyW/lgTmJiOAZmExUJEYpOFn1PZXW+Ioy8e
PhiPL3oAxeD0EUbQIM4kFqBGwRDK+iCx2h0rIFZi4in4+CmpxFhzki2dGlowAzikN2t0fYJz6+Oy
X9RtO7jjhmgtXOndJ05Ajj/Q6Rq6Jn+lkVPc3LqpJQmsOSPhXc+hPnd+5YxWPsOIlgeEzarzNhZI
hyIUuWHPomDRPk3llmhTUD8BHgGzHONH8xqD39Hz7R5yK9Tmo5O3thFaFUs4BtRTdi1dbouYy5XG
c4FlzA2UhIzYcg3Ds7UM/dJ3ywsOnd5LoS8BG0J5XJRjgBYkzHLbYS3V68hVMgpn1MEdubj9AdMu
uaxv/E5qp7UBfg0ZiXk6nAw8Mj/EFzKrXczTJFFKBKr3MmW4QdQLPscZmtMvomWXjSN+HLCDNojW
e/iQEixrS91eQmDrwe1V5xFAi/ys97CFUgE673CaEH12PZXly55DfHx9Rpy6INcp3TvS3kUE/H/v
4lK09qjYQqccD4ctBXSzDW0jV62SCCDWd53mWtfZXCdHBoZTUHMaQppxFl5IavO64xt98017ESSL
Ih2ww5XorB5uEy8IBwXpQ2s9BcUgaRWJ/zoWJlTJbLwZgObobX2UyJOlOu7KeIOV22iwq0bZpDfk
mIPsOfaMqIAyBozsCcmmOEHa+/8Gvq0pPaay8VAxbGjjJwOkDEhTOi/lzgqKu9DbvgFWyZm1QRcs
SmdFfqJh9IRu3dq39bvTZ6HehMyjKH3nPVJbYmEzqyr1VNIcvDBO9B+/ZinVOGh8OoDOWH3iKyum
i4hTomAb03YLKv69m7aDzzRDq8Xe89KZi+9D6mXs1siAYP1xCyXN5dicTHoPcpGLeNTGkwq1zjlU
hKVM2Oyl7M6o/N1x32lH6jejpOt1hvrWWmDOX2rP0K/8vLpVFtQxF+9Q23CUMl3gX/hVJJu4uqMV
7WAKroj7IUG/etstYgsxnBVgVXUkB1DMEnZqiCCVZhI9wtdEEPuCs9xqxj0OQRAmJ1i19QRXXjoz
9Jb68l/8/BxaG7jsmv6EmttOucE69OBLGW2sumF5S3agtgwptbQRnsxbDTIH5vpY47gw7o0ugJid
m4RBOvuoahfJLmikvCeo7vntzh7eODvEoBt8gf6cB1Km7Hkr0NkduJp9WsNcm/s2t0nOO9alf7Dc
BYHNc8hquXrzEQAf9160mQnlOoJcWpDQM33QHqOOADZH9fLszFSPPJtrguFZhCQnEQ96XVo6ZFD9
ReUvVD2FM9eaI4bfrSPYPz2l9aqA9ZWM87DfQlIAT+is9kd+HOdn3uRaUdX6ocDfLSNdbqx0kVBW
az3oRh1ATTMqJpJ8K9vqVJwMlGYPVqX1RtOoKMp8udsh7gK+axSfX91Z/315AYaC3qdpdxS7Ea0u
mjsrGwOozK3nJY01qv0x+2HcAxH95eGu4pyPGRm6f5imYlVDO2gxaxLV5ZYFH4FAYXRXMYDPDbwx
BaiEb6NvMwsiV4qvpqUeQGphGcdgfdpI0dfPBQ/QgwfBNJrhC9ocPlOsA0bVhcGd3wgzgP7a9iEI
uzt/Hp+s+EYjEj08CvHkMi/69j4J2ddJkrCzX7Qu+UWDlIA+W5IF9zc3XT//6pD7XOsqn4Yh+L2N
1M4SncWJ/kVswKSLHIxvLO8DGJiY33JNS14q4W28Z7dWw9Be/vG7ZWN2O4JeJhuXsuzjmsJKq9fS
29XYKLxHVSUNqIFeGJKAtMpS3p/7aZ+rEqLFOLWy5z9uy4hgAvpXrSe7xNgugTNavhdn+2KKAvEr
7EhJg9zGPnT6eG63Tsdi7Bgvf3mBNThpim3I1sXEjozwqmSZRg1/kt6kiOkLvtkJLySv8kHbYLqd
hd5zYp5/6/dO6q6jseIlq1ApVox/m7PdxMY6RzTRd6gBV0IWJGzq9FU1AO+/4ZPfmxea0t7KXESf
IPzgS+gTHBQtPACXBDgsOIjMW3afZOhmorzr5EkST8nrIb6sEACvE6wPRPklYw40z1fTMoAa+L6C
BLita9N/GoM9WoLerJ9xxGCroNfRxBaZtiazpvWlrmMqLWUuRwWynnAQiXTCrqPcZEyU6jmsmrYb
coYsEQszfPdLRgRkuqAQg/c4RNaDJwV10T+4OfKHTZR2VwIcxZO+K7sDwxvwkbPC99oCz855xLSE
QmPbj2yqkrS29KG7lVRIfOV1OOwoS5+k8Jl7bQ33iawsCp5jWNKQzN0MsMsfdMXb8engjXqBizYE
vLHGaahhiH9LwQVRYWKe7xj9Yjh1GQXG0BkJ01UMr0+Ff/Y2BlN/hX33LpGkXDP/KOd9MIbW5WTc
S3RgpDdU4hVw/oNA9PbXbXKhASBN0TtObBeh7GKOrSiP3DsYNj8h8rUukbmCH4+hjz9JQxrVE1Df
1k+Yw56bwJ5pF5nj8q4z491wuKVjBFKuxparzR/xXKrT2NnAF8uTgC834qvR0cDbWLw5YQa5+9CX
rmC3H3xc9qc+9XNBD1xoLKqbC0FZf2kU5s84l4ybXlcFmhnlqxaweNDCzSYuixOyW07zwD3f25EE
9b9OXXzXkaRjewIziAblpsNw29JieH+Y8ZsXa5XkIlC7c8Or1D64mv0RmphfRlqLWUBMGkhYhI15
brxnf4B9boiGb0vs/d78/Td9GxxMBICR71uH4oTbbSkbUmqJc+jHID8gtDwxS2Ft69aisccmbQVg
d9kOBETyXTsAgkKV/x47XE7im7+pkFoV0RugY8Azg1SL/Pt5lynIR4mw8PpWVn1R72DULpGLvI6C
AaHG2jXgeD/lzhxQEFinuyOzE3tYVQP+Ft74rGy4N7a/d51BF+HLDij97GAJZsJeASqjxYzzFavW
g4TgzJ0j+iRSOcszQwx8io7KcYOT5Wk3CZfCkeca5zwvSv4epWd/Uikwoo/miqQIkitnoC25Iomh
Tvfa/uW0p4tjCZZO6yiAUsUeTO8U40UkkvD6npKJF/hcV9wmTJZAVvSG9HF8tVMycuxVCHsifaBc
kbUApgPy3MImuQq0bqUgUQvUZkwJi7IeBRnhliyZrxipcSPnbafiCUqYZ2hBF2+XwU4+oAM3C/UD
DOMNB7aCyyB/08Tc36Pf78F+KPMAxZVW1gVGF/vI8hSiFeTHobkKni682Jigdaf6WUnJnqtAIrUs
Gd6O9qCs9GHndZI0lxSaeBxMb+DGIU4qiHwBl4WjgeOkBrGQkclXVg+XLeRHTIllzSYhiXAhfA9t
YbJQkFGYNnyDNiyAsgUqoBab48ecy7ObAsuwkKN+GPc12rEm8A0hvVhLNUBz0IdFTfc7DGkWYsGx
UEEvcIUVOEtAt9ZQqaR4HfqwjvYkCjS9FfLfG0XJUZmj+PYAkBJs7Y5juFC5Z95amepOeGnJy1OB
0tj/70m30zv1r6KOz6DaDDY6X+szGw7r+mc+QfPlYY+FfPxsr0W6kwGzPlpSHKPIcNZcuSZzZSYf
16Nk3+lHpk3+tDWRuMe7N23fEjXHXS1SkIqstxsDqp7kE60blIpQjaz91X7cjjdAv8tUfvkB4YHW
xTZIT54mM2b2rVkOW8JOydCKesKIBpqtCCTMJQs0Kz96DxRA3jl3X4cCPMDE0G3KctCNkTXQrgQd
FyQHjaSXbIr94CPI2xxyXtP38eXiiKyVp8/E3tFW05KW/Ze5ULLItw7nYp1VcFH5mrbHyqDUMy0A
f3QLr24HRZPpqHG3Xn0lu4KBAB2ZVsf+ZPDBr2BJvM9NpEYAwzljkx2ivHif57Jm79x0Svjflics
UFEGoP9GM2EEAhZOn+KV9B1wPtUqZgV2UwGn7kr6baiOcTC6XuluR1VFvmmKmOIGxxSwna40xk/i
npdGfPE90EEupwYvQK1IuITwFdCknWlj+R9Hl2V8CgvqLUpM5B7GVGQdBq07CfCaaivAA2yvt2qf
I265uuacM7tn0gvAiTvKYi5xQ7JrbeYrByNXbLNO+JC6i0VAH5C93At031pxwnzxtn0+40w5YIwm
rn/MSmVpd8JSTV0DBFughp+OfVmZ3QCn4cJqgFlwdJDS7Vno07nr+ds5VjKTEx+4X/mvnU1J5++R
4g32i51zNun7kozqBmn7SGWG3x2zP2ALxkzvI7T9AnxwCxaR+sC/q96bTKmoSzeNLARLto8ZCD0r
WkEIQyc2N8eXUZDBofahGTwRI5LENoebUo8Tev+h24YuFib3yYL4uxVYmskjKTm6qzpkMUIDSxaT
P1gRgkWqneX7SPYJIes1bgVvTrjDf1Ag5Uoam2uDAI5ZVoFEQ7iT2VSUHmiGygPZQ9kujMknqXum
/7rl2ZEyzg3r20NbkwIwTqbbHqjTahINIBPEZklQPodFrYGrbEU43rFE+6lR017P/eiBozod6Pra
SylU2roralKnYEe1YyW1q8+mfOnMPl8QLFqCm/4nafi5vFvWyudsnY7C1DjYCXSQurjeTr5Zci59
tDM0Z1TFmWg/EOjzcUFo/kkB9lCPzuIPbSBZFiPr6308RKQo/fWdxD9Os59kNXtPfiHTcSEXQC3E
Ic2qAQ/Pl3q1ELG8+paovXxgSbxDbcm3LC/ToQB/OUPUe5cdyWFqSjQSdY22X0+se3JdNpQWFkqr
dp77zlkK2Y29HAFJJ1bsDmGOZRkUR0k6Z/Jz9dYUnXZWbk3fhd4cOlk/MCwp+8R8JZwDnherXxwa
jPbFm68Ws5XuJScVmMVQYcMV8P9cTpXlX2Z65Bu8U5FH9wTEXn52zaD6f7z/9U4gsYXWcrKYROSF
u3cECgTI3rsoLhxesxjkg3lTnhpaBjlF/PJWI1P9MVJj3xNBIwcIw3kMzc01/Q1A6sOfBbtwVhKi
6FmhrNe4CuzAM/a8gIdu/m7cfmTxttPs0Qk+1HbFs8KRGLroysmEGJsq6Ar7Ai+Jv/DT3EKIkSLN
KC8Lcqr52L3i9h+bwWT19JoPbOnATow45YuxA2h0FRt0za2KtvdowHMYceO7CbVB7dXzxfakxR+x
khFXUyPYqUmmBKC0pKwuc/5qT5ElZa8MrYgCeFA7BjnDwxM/2+7lRgkMJUk+cjg5Gob6YBYqW0/u
KlF9NJQ5zOlVzetjmDNYxNTRA3mcBgVwiB90yQZfQeFRBwLvSxBQPtzgoCszMmnEcnmx/blF6bFS
yp2wBJgl4XR9dJNobJW9BMoDbbuB61InZ055Nht7/5VhkZRTPcj+XRl4dt1w5o2SvNRn+TEBWvrU
YVBXM/ZYcITwAO695KZWnD/sQPCWrQ3XCzte7BlwOxQ+kee+8ljzkFophpFKiXkq8kBjP8kE4WCu
fUTPI9E4Hec4siOyUinStbkaIZCnA4DDt0K/K5dWgIDlc37phwq2dKto4KCQI7CzXp45MoCNfTpp
r+UzgFCiIlBqiuUIId4CYWAG2uQtX6k+CgJNz6L42JJj2dwrZOMoJGDvusQ4q/8HCr1krUuy4QZB
uyf1C9dMZw4aEXPU3wXC7bJnvc5gks4HiGO2rURrljB4ZUDvRgH1MQPnLR+RURqq438aa891d0VR
Gev7FEQQtBE9HVkFioXfpKTp4FtOKE0Q9Ukl7r2YQSOIuiglfkz4ajXVmzrIJXHRbqFirAjmz2jb
32CzNaYLfy6BrhFDSm9o4DOt3pK5XC9Po/L3erJ9ZKVhhWiZLvLgpd7bZ9umQtW9Hr7FvGcCkGv3
M1NoqG78qNwqXlDWPkjN0tECCzOBkBaIF1vrz7U0vNx7LlrD+/v3BgcFjtj+ELzlGsDolTqqfC/d
qQjPQZ+BiUldoy/t4NzBerjiCVt92RFaFLxiXAtsdfJwWqVCIMMeNmS3lIkEeDVq2dZPh3ZT9l71
mOJoIevcob+uawO4f5rA3y1JBVhdSHzfzmbG3HmnrLTF7ku5UzQ/O5df+mpCEdrqEvNmVbKTYiK5
aN5KgXtq6I109ov5AdJ+TyvTDJeMaZhoGLRgAbS95ybj9UwFLWVIUqi2WkgcdTEcZVe1kmf3SBlS
VyR5ttUZ1boUAROjBdzlv8wWKG3VTjXoal9a/xtitAhHellQ4mUzypdBcODNFqp17DNx0CED9YtS
1IvRQXAI7qgbH1uA1Gp8K57U7hYu40I+V71muaJFlApKQJMyXPcBqlufOmDBIuLpkYj/0p1/MKHK
y7/5drN0Bdx7gfjbifhz+a0Q6WtUU0awQnJyWb9GvtuaC7reN3PmCisT/41GhfGvJHjbEGwiIYKJ
VGr+m2exmkTVqdWCabdVsk8Y+WbDukBmbi8lBpsylFaWnLvdpA8ezFncn7uDqHZYsZvgPCJ3gpE4
usUSlv/6xtgSW8HrFoF5fnaFOAqrXRCa6ijfkWxNiXc0cyMpzX1r6dDxU6eTQAWXZ2I/P65on1GC
EuxqCyqDJJaaCF7P2qSe7vnUCkVUPZdHe2tTZXD+2J9kmdgqxFUa3Gl4nmCi5VuTtfJHAU0mf3WM
sUFdcGTgZbWv+8pfEWqcIEAT9RyyTs1VCIEvhvbw8fJKfg6cxZonQX0JWcLbeUlyPUgpneW70ofk
1xnUaOhi3CncTvMhyixKB3e9ZcLyzdCCkmV67TQk5tV/QYuMGtEhDsEtn6XiPpBopmg6eCcvs3gZ
CjazlffkyClKNUiuCAe9Jurb3LXqtZfDlws1lLScvGN4fSC098f3H/tz4bVwbz6WUPnzC3pJPEKL
g5c6iegEL0R8v2SQ72KzVF6zWz0Ypg4kiKiF7cMO5LfjWtxhrZ5EyPxPmxcZB7gqQsZtkx21e8Q+
F0OkuDo1pmcW+/hZFfmlKfDpHToKRF7sf3u3bBQCSnL8BFRQggbO0OaYaOoQV9exDLCJViaR+Z7L
Shjywd++yKEMjPchnMT8FuHHjHpFlKHHsd9MLCBXj4MDZYPTXKbajWKv6sOo+GY82V/l/moAifg+
oF7vdsPZzXa1V+r8rKKeM3tknr58QPYu+dZhzOH3k1d1cIA7WJDXp3D2o++24r/meLL6I2GyXglA
X1QO5jrN070VJmiLDP2Il5I3lWmAdUA//pbhPeCpK9zy92DN/sE7KNd1SOcxm7hbmnmaWUWXQ5r6
GnxLReX6pp9Eg2CgOZAv47AHEBxNidPb0cCGQNzsVkTmAXclDwEye3pEmvLHgP8ZWTnYqiy8+DqP
ROKN5IYU8iugx9Yn8zEiewvIjwXIouQBnFm4h04xW3hWQQ3KGwZa7+JB6ts38wX4KPeRIgRtbmN+
sPg72wAABzMzE+kmdBAxPCq3nuERcm6BN3CxbUvbDhwQm+1xJ6B7OX6mNnADErdx6zDJNKPDtq79
HQPm+rx69KKoiSrrgMv4xdinvC+rWx9T3qfDYvWkAqrHJ49Z9d3hFzpk2cgJ4y80wX5QUa6PIned
nPTbD6ITYrSPi6RVdyPsUbW9Kjlkucx+NBQS+lVsjLgePzEg1hveqUKIA8UMtNqhhqDLZLVj2dtg
Vk5tlwPam1eD0TcC48pTvtZHn/RtJZKQrxdPvO9oQlg+A1YDXhrkclE3KM4UC7EuZPAvuyDV/c1v
IWo401jxfhvI7epOKhSuNC1zBGZpkiztVNcEEQ3TP1zikmITWAOgRCuTBdUxX+4IzPpzDO/gxgCP
WoCJnahe3hjxcnO5C96WHZi7ROC8a/YwMhs2Z+nvCqNQo7DZ5eSc/OwNOHBO1MavzbjTe3H5O5gL
RrLj5XkcgZ40cQgwa7YH6BLGHPq7dI/lJ+Br2g9Swkl9ejkpxT6RpQE4jBZKzrpXP3v+HykTeChd
I4X9pej+VLR9zwX5jjQxd3iZJaN78Eo2qw2gccN+9iw9UT3qi9ZQ5olX7YVpmzxuJRtDe0Uzcd3e
8LdOHXId3ryNVINFT9SBkuQZPME30xTtYzTSCz44HF70vItQMNh7YtD8hMmQvBZjfWjZwPPLfJ4T
jXVUlvV2WCqKy91BJFS/PEFjv3yJLEtipR7WsXfpVYRN8rxrPhoIcvreIVEiichDGzuNVEhPukAf
8O7PltoaKzC3KDlSrZkRYydfWB/IaCKV3KzDqQlArmbdAaq8gG1a5i9VfQBGKRRV/aLai10g/Lta
BqNoNgBCIGlhPy8ou9sOX2BD1WQDNnjtpeS+Pm+Cr34kz8XXP6d6KSQHvxKDuTIlcXhE/5fzRA9W
quL1bM/O8dfEpOecbuYzHjEUVEoHehtGHq1n0TtyaWOM2r/KYJA/mxCyCUkxGIeDpQmaVMSpqSAx
q9nHRIV9GEke8TV1rVblWtyhc6zxnkP2W9nK3p11o4hPiFdR7YnRiIay/d04eDIEp+Ipy5/TEY18
KpqevEHtjaYxdZMypxQ83gI9oLyGxNsZoww0mvtpWMrC29+Bnx3IejK8M20JjYdZn0KVvv/YggwI
3wYgUYHyGBnH+GUUCqKmYmA6habG12+hbmxsOu+5GpVYdckjlFzEswKRfVj1vxjTo8bVBWoeiVZ/
Rz51r47vlO8XfyCefvjCx3t6//anp0gxp4iCiHJvV2Sls9pIVR0sfArsRzkjghYGG14Sr8lA24oS
kfBLxQxfZncsZ9LrM3Wxy+LRXreDZgJC0z0PipkMbFTlQxwmN+pom+rKamqgyfzG8QtEHLXGdk5B
P4A2JcMQJeQ5V61PJM98YZHUY7whaOiniXYdmb8gggFy/BbiZKQWDvG1xjOuijx+s4H7fxtojKpw
QJuyyHHAhGuHX+PeJZ6gTRaxyhKivJfVo0gxxT44Zs6ulMp6e7T519P9Xa5OntxczRVtub34Md7M
fc89WuPQ3QLjGCTvXXbVXl5cF6NDhEFaO9HFKYRf9vs9ZYduA/IKTcH99sGmYc77/arNrhAI1Csh
0jXzi1uh9h4+HdE91hAspnoO4GxU2HHvtiCimirGzstlftRh2dfsiWs8mF/jw8OcUKrR11jA8VYK
xqX62+naaYljNHwYEgY6w7KvixvkxNH6JQtCdq1RbFjyh7b3UM5eVsR29DGMtkMCpF7iU0uBWGdZ
udPqMP0uhQ4yTcjXI/w9bahZJISD2GtJ1zQnS3+ZIfNSgRaugBtz+XKqnImo8mpFefroh2Zu+gKq
zrzXU7sNQTfDqxMAe17R254B/YHhTkBbFNJNXJpCWi1S6ceBqDJMKaUd39pEqYya00KQ8ilI4l02
MeiWFgJym3xVAlZOIo5lZkY4JzlK5aE+Lwo4KV4AT1cXtNJRsrTuadRwv07aYY+A13V2Q/IL5JQ7
AW5cchXMKr8TKfC8qfJgMXmLQvl5HtJf7YGJ/AHLoPGL0QPXLKj6kfYTq946oxstYqk7DrB6ct06
N0xCc3e6WllIkQp9fMhooeaC/5tTeIU1B5TVDT67YED2r6fpRp70v8fxtM1pHPSGUbEpQd9ZpQgI
D/wniZboy6TmFuJttrLHrZZ3xLWjxqNzyfFK8twfnxQ9PAwhbh7HouA0xjaVTSTIlaSrucDon8gO
o1cjPRmbGvO61fXKiYN1TEwV9pSzeHjltiqjGBkAVeFPt9wMgZYyxjMMZbuny7uZgDYBArFAPLJ3
JoPA45rVFge68K8XNUyDsO/Dv1V3koR0rL1gLXNpdHg7ehc3CfANh1p3JcTxkOBF71xQR58SMukS
sucLYYMEvKQHBx81wjRxN0G3WWlFj9TH9ZyAKhvbol3+c0mbo7pafHfnjuwOJ+ssSOzIrE9nXYZk
J2P8sL8wQQgjI1jAl4ZufbVsE6ngQEMDiaVYwNX6CFekH36B1b128w6GRXVcvHgj7rZCP2wJz9Zn
uWR0dEMTTQu5X/oh8DglYwf0h5OMvuuW5nGsHaKuquYmKo9doiJzFp/UFr8efmGsN4xVwhvLbTPn
ay/EHuDDVNC76amgUmGDsKU3wTcuM6XPZ7wsM0PfEdgG7FwLmvCo3q8wflA29Tk51VEGgHrtaKF8
VHeGDoarfh/VeqMiO8mtfYUdSsS7PSAo0Qtfzp8yZ9BLJ40NKSHNN/3ue/5tAhgMAEKnVkA+Tujr
8gQB0+TblgSVVMqVjswmMz5C5nzFs91Y0maMr+iACyuCoZpGdzppnF8O3YsRkj0oPhSXMcdHAdyW
fwFgpN6Hb1vs+M5ZcRSaNhlxc7wxLONxtSRvdqCXpLhEounjejdsyVjJdZ6UDYc/LZXCErtJwM++
bKClxH5TCAGRS/F092BiiX4084cTq3rI97wmMe4WYyBsB3i1U5fzijPabeULMXa29hOQ3RcVuANA
MI/diZa1ZPsXFmVGi5L0sg6DiEY/pdZPpqWR4V1DBrxAwrZiXxr44zacrL7RpfxCdyHQAX6TmwLy
89MK57ML+BDClEaQwkONfEl6yTtUaSDc0D6FrEK0oUlG60j2mU8NNKp0oJwmND80nGGDR0SwjRiQ
qQch5h5sdSPY2sW2M8GOE2Xx3E82VCG9I2lDwkP9/84sxY1WluidO+YGtB1ThXpl2m81rUh8sdjE
KrqUwBW3Bhu33cKEJ9cyBXKpOewaGrOQ20lSx1K9lXWWHFyjRK+3Xaf64sUD4oC/HQqA5jmGUUpN
jGHvZGLjXhk2uxYldmE7AW8tShXCQkp4Ep6BxlBHhZ9hD0ZC1X7D4UQHSBwdH6/M3fWIVdSghSOR
0xuQHe6tRbzKPzQdGSQXtdZFMMuFptGsryo9cErFhxZllZFbg+BE169R1q2M1I+niZ9lTqpY8wnO
2iH7vV3c+1Izv9zG53A7BmG/IQHZCWyY0uA+3dqp3ofTZeIwZ/cG5kzp3t+2fq0WmGHiLX/EQShz
KyEI5zBkcGG1vzwaAURqtLNeDVihPtuR1YAUdPYRwSydugHWV6vquNk+nukVs50+AJwthe+4lXp+
upcBOPNads/xqFQARu1PXNZrLozWyz3O0e4y+Q455WVPisINNRtDTgQoTadZQREzdTCnF3j2zTo8
+CbMaC29A75eATxshZGE5Aaqh1+MlvtVwuk1TEe4h0sitbImmPFapSbr9RFvtY979TDbWZu03Lsq
lu6WjH4aMXNvOvfo6LvMopX63W+9k74fVcbfFaoJcnpmJvKwQSYwN66auJWL0w1gWcVsW/Iuq0WX
LrlU1CZ8vCNE1BbzzO7RulEaL6+a31E/ytj0cVQegCjjDu7stN66EAGwpG15YMU3xDgII/eJmI/J
XGZuhwWZYOgjmUdgSu/nl/aHMDzjMo4t8uIxK5ftwSCyTgFq5g0z4G4QhnNqQHMzHGQgunzrXki2
jhVMU1Q957k8It5rAb7QVrTtARba+Fnvp6Ad8Q5uQjLd6arhlx7D84k8Ylfay/RqRNmedXwx+tgE
rrLYfyq5XZoMJVIun6zRBMj5LOi3KQY2ILWyzXFs6E9nf5tk+zhuP9vqtI46h17pVjqYyKpvfPuV
vXdgf2kVEzl16dr6OXTCwaMPUfx6fD80c1YPBM6KkGeDGIHM25ji5w4caer6ZaQKmlA0bRchncQQ
wbpchgEPmCFZn6qoak9TbfOFp/72Zo6KgbvIqyPfD0Ce9XWRs4hQsV70i+gg0nglMd+dxSvcfT4Y
t21bdDVhQG1CwuhIHaXioti13g1dah/63RqDYkneOqzlfy9hsOuWXFdsVJj4CIp6TfPnC8dm5AeU
ARUGHw97AcLvX56jWpgocc/GkZQ8ZuiGM19uTn6UfX3vCHCk403BFo4T93N72drhZvEicLs52ufq
/KXqp8AgwS9k0ZygjgjtTFnojwjgYV5rmNsHbeXwMM4kBXmg46OQQiJe8wYR5lnKPlLwHdC1RG90
zC7cqaPLyHe8dW6KjqH5fGAu1SevHJYJ/kwSu+52qjm77EgSLNJyl5OaB+tZKY0yfMVQmYcf7tvH
IawiGXqsKRK+tgGgKx+dMIy/FA4401JWx15B3qbb6Sf51CmHD6wS1Zj3vZ+vpj4ov+j+7I0QtFel
WfYglWAoYjqtt1EWdntmBQSD1/r970fhB0T1zPBlUhGDvSc7I3Xh2xsFToZoAH6Vyy5TKJTdXtnM
G24NDYFkaTS7wiFuHFfftloOx4n8smFb3g/jcjbJ5zqwL72jF4jt7SzQPJPiGE53rNtubH6Fkgtv
IGTl5+C4ppwSUV6xqX4TP59e12dfOe1YIeX6UQc/6T2kbjUjVBhobguZvGm9UJuHrpZJImuO6YQd
gUoZGwQK0D55MD7ojxpVrEGoVbTmoeeDTPIeGFEHQ2ZIUPZVTT3CcqxbGJNR7hPc6P+X3wg69kcT
arnGqFh5TKfzybX+Etz0pxGhW9gchQtsHXCqAtIPqYyRI944p5vbqlhd8cy6ATyhjbKegsioNT/J
yEz3sMDQdmSEAHp/3dq/9FZo2fGY8jeOk3u7aNUWD8Dxc9Cu6mNY91LUdHLjnC79gyydEFy1W5dz
4MJivu9Lugjs4DOzWGot4fcqLJznakjzUu8vN7W6+/CNddIOJSVrOFvhTDFQyvGk1r4qHFVkr4F0
PgmWweoNyyjFdS/yI1mk/3OPIKXwZxWGk5niVMTMfmdXdyKlDtewG0kKvCESMR/HD55wcAV0qaFT
+TeGKX26VCs5hP7uDzjxIY32YmiBjdCKVD0ArpYlagYXp5PSOK7WhKJuNvkwuyW11R8NHvttSkqQ
jIk1PmmLUb6lgRbtWvwmcJwCSNs/OpDJhpwmA9Mwty/riHH++daGyNueniKjiBM5KIRdLMnKOxUf
+jKHmipBmdfaDj+ILSjDowLscx1zJGjLNcirWwoSvB0L5teYIX8GK32xtXqjMVndIF6ZYX/93UMY
dsmayrjsp+BqG/AOzu76fFx1CQHStRZ5cs3Mjw24HrwjF8o8LbzSEilEjgCZ3bLnruvahT9Utc23
/cdGvmpg0g7cXm5rwIPfgQhgfXSa0jLPpbkrL0GPFhOsZQWQ3gq8sqQSCmNmKvUUUxVIcF5x1Ugi
Hz3KJnBV6JR6EMCDobVPo91IEZeWN2DDfOWfO5yGQDJdRqhebdNq4ylru1yUi4zUJK8/3I2NY+A9
y5iTR63SccNGIgTGmxhH/eXJgG2iDGAAhuT08t4AwPzSmGq2uE8qvZTqU5aqrk+Dsf+1XU7Pzm3T
Xo7CdyhPhzEHp62asBLAW5wolUTE2VM8sYmxxvdzenmv/VIlR7Gr2Y+8uKRCWa/CmIYiTLOJHMTW
UxWIrMTNEFfdbKILVW4DsTbAx4pjvYAReHwgLLKNjwBooVFmMta66Hlcu9jsdttcLUezKBYBaKLq
ymSHPJ+rcRs49EkqaKjzAgPhikNhALM+MgopHlprPhrY7Sx+xQArOG84RY8MvlBVGdmFrOQJJaGa
mwT5sti1LwqNTlYFffa9EMSKayIKU85NOuv0k/9gcf9hid0BfquaJE1V+H+KYPNWoT63yiXUEBg7
7QVhwCRUs0SnEQhJHrNMy27aKaEYqVNX9kvW6sZbEwtYdM9PYPD3XvKeT/LxeU4TS33UEGInPcUc
UauwupW+EeUFh7j2zBGnDevrp2H1z66e17ijEp+KUM50rc3f0shOKd0gkYRnMVHNExaftVInBC5q
PactbdOpXnI0fm/Nb9DNrtGIJWGGu/WBjMIY8hOABeDenFTHbdtp1YhTRRHlx7GT/+WWZZMOOvcI
f15WJ4zl4vUSQ0yNcYc1/83tEw/qIybBYpqwISsNiBXfxG53pkzyHyqE5q3jIe1enz9S3UyY1l9u
IJgEoU81vJU9GZqUhK1hInrRtYjX2HGXJ8w9YJ6ns6R9fXAcwY7deSlmGpd9m0f96X/Nb9Bbn9VY
WNRq7d5GjY+47MvE2ZcclVRiz+1KPLIqy21LbL51mdP5CreuWji5fnxeGdnOcAQ+qXB/kfHVLn98
1zGrhPl2yuwZ4XfBjq2gVGWhPj7sc4bFzQ4B+XHawmRIE1MmxPvSE48iH/e7ZYB6/qnyFk8sSMwF
0cHZ3gLsqt24yFQimwEWdxthxDGbj/7ZBakmXLQyT8uVfBwqy0s9vm4mSEpcshvb8xbyFMhCZKv/
xZKq9D9pum4YghkzQqboVXf2ArvHcAu9gwXDJr/iFgY/sfnwc3DOGPyB+vHy7Y09XV3GuuCwqP2R
OTSE4L8Kul9xcjVi1AsyX9QZUPKxAybRf91Kwm1Q0AoCEjTDkvvqPUsTROdIdy+ZUisiYffKNlvh
U952ejJlmYnPYdSp8mpIy6mUh/aDhEHdMuecGHxlNIpjgRERbueEEL3CbcVVm3F2zv5Lau5rJble
SQzK+YQlIpYOsccuuQ6u9N+YfCVmFANh7GPMTjo3pI0kX4F2LKECTwi0/fORAHnQh1NNfQJjmknm
wy3F+zOlLRLb4Nm/L4mDt1K2FMif0Djnvsij3Gphgx1oh3KukW0X+deW9W8U5D4Pxnx/VsXg8km9
wBSjtw8uRAyj5ESOF94WLDhj9TsYUz6Y7YEcXg+9zF8+b24k/w1d3ky1kZCHZfBZcDWJxyIBThw3
o52ua0/Fv5S2To30SXDxQQGfmzs/6ojFq/amW3odJZkAQuYUEaan5ZsUSqktwq4kyE25sU/iQPQy
OaNVuAEm6LellQfkWmMwBHu07vOAH2QMQozt69J65cIPi8Ql5RwUFpx+v802Wdi0Z3CdMwgvje+0
b3fED7PP+mMzaDzAyNv9XdzOlZRUaJto+1yu1WIIz5VycsHFmE+hCMh3Y4LhquZJPx2HsKe4ISd7
2ao5/1nk+uxMUbpz/C5hDZ/DSWHSvzL2A2Bxprl8lwcmResw5tI+fdmKBwde8Hb2/2TS1XNbT3gA
9XDFj/tl4B22nQtI7C916NSHMytk+WPP9nxTRSeL3cn7/SilNdq88oSi1y0cazwcUgvkBOW+UDY2
SdAyImPex9JCC7TQKqlaDv7bvTvJHQYXQymlnSW3rIWSdDFQgx6wyYSOq9gJXg61mfkIWJV8/kh3
81dE4GWnRmXmEyXAiy12sq+DtSQm9Hu9XYPuHKgAtAsnThjcis0BquSX6mCTIs96/dguqfXgM7Uh
UUuolJn4HE8TLUUnCLd3mJ0D1lC799w1oZ+P6867Wifgma9ATjuAOosylToQhx4jBaCG5RG4gMx1
ApAfMl3QiZoM7/CvexoXsaLFoMyrtLW0q0E65Ns9gz41LHP/H+PXeG7CXz31NM+xQUDL2uhTaWWq
2fDpypvaqqOXqiC8ivKxnLRA8WrCGaSWJWSTIRyeEcbEnT8tV+P20cErr0vHqeiy21WRBgyxhEsX
q7Zd2fnPpcX+VR2wY8PPieE91/W9xqQZ9WLFmBdwMynDDXhDteRHXlIVyomeKHBd2lw0XP/VSS83
PZMjqXAQlJNfoClsIgyRSd7FyKtmmC5MBmSlwHEAVGkmP8Oh6QDwlSjz+59Wty9OEk8v1pyWfZer
BA/4fei+S2HllWldwgxPoiG94yZRFYBiVIBI+fsc27UeAUUnrQRgyZSfi6FOy5aTW0cla+9irSkh
QMIrHbUynXNo+3BQf2M+nNDB0ySEwzcFDKAnAF8JF5Rh3rG4yS9Kf4BkZ2GORACm5FGmEf0umdU7
zNY0QKNkmH5NGzqwEeYTfvIdWLbUeelgkaAxCMia0FeAp8EGwTtHSCvjElBmqJ8fPlvnaIhaDvAW
RWXWSOLxYS8BFTz1FFoP9tPThvJ961VN0SblLIiKkCbjoKJxRR/Pn6oz4ZcAU1LRFIpEtIsiax56
8/3flU5KGeIUn0sZNsnaVPevBPnaxixwrPY9U8EcCpjs67hJQ8rqgzvNx/AHEQalPXKzC4lFrW3G
29J74Oa0AN1CVn7CzuSkrlwJNEfJPo2457rGOwgZEfaE/wHKPi4K7U3s1QuPXZeWn2Hl4IX0xTVZ
VtLxplutl3YtdliBBCE6npZPrxJZzu+Z0qGYXUtKRoVwe72Y6M8Fx4xV+k/GBQd83XpwKVyXCyLO
7Z8esvdcq3FH6WiXTSdyjCzdwYqRNztQQj3pKl2rj6i3YAaId+uN4+elrJW8RWkISvH2bVDC0GV5
nUuQ86Gjs6Db9HDN6ghlxTJDrUfYynjMQlJKF2L48dw0qiDtNa2r6GrSBaY5pBTXS/0e1BY1TwoW
pni3sORgVSQ07ALkdd3/FJXaHx3wkgjf/UXTliQtjZBWcg/JYLghniF1uw0KE+WvUV1BkkMb6vcZ
gVIpugvzwazCkHcRhBrIkvSufeMr03YMUsAfjt9RbzRIw4s8vr07GgjUJTLDJLwhNilCj544iGWX
MG8Ka6c5pOmbyEAOuWW24dsN0XysTh1WfkuAbVvckC+l2uCNjFQTcSk/TWJPpa3r3q1HHnmTm0gs
cNn8x6crFmU7RwVfBeD0NwaTFk5p65nZ5ElIBCmc9ll4bWbdC/0zeeiUTCzGvsMgY/RXKrxcUWJ2
P8CsgqX9sccvnCMZV0syOypO7PAaW3LkIGgie4emhwxNb3jB3A2xtyuuf7R6ZUc4MEX3aZTrwF38
7CdLiOx1z5HTa9ZoBB57pqrEdFivi/bZdFMbVDGFNWNJEOxEsNcOkT1SFFiMMRQrLOz4IaeSwzIE
+5XXdoz+Briye1IP4SxW9HKYcclDGOOYeevnxgK2ttomKS+YM0KnduuXtDUrJGjMv1IjBrraeujn
GD2IBz/DGQiLnsz3QuChVx87+UfsOS4C5Q6aQJro4n1lLlRQ/4LhW7BYjMDWyOspMK+yaQJvY9PD
748XyhAessA++pHTuYbHpJUzl28iXgycCS4AC/qy7LLaRl0H3iNpUtbnRLh9nq/HzCAFS4Y+601B
MAjAOruJqGm310CdNb+PbHYWv5GKGx7bKNkSz6pHlsxSeTXA39Ahsu9l0PHDjqAj3t3ymN52qltS
GGKgIzYAN1hycQMNafFND2Gr/vt6sh/SKWrX3rqV1BNJNF7BPNdPv/ALnWzKVcx/T5OMseU+C4SZ
TzHA89WQn9cFjIDmFxStkL2XacWVynYOpvl30C4kYN48U2quxOpmrpJ06O6RO1sMNttqCUAC1/1Z
GyBKco+AJocoHj8Wo9yuKXM5p+UGIfF9Ir3t4suAphZgy4S9Pz9FviJZeJk1KjYhTwnbIQ0T9sRA
jZmwHv0RzDZrjo/J4IcmyBz97jYUbpH5/PHzrXr9LqhYZBLEqUrKoAqQUrRNvqSZoBmMk5YhLl4e
pZyP7bxxz5b+bhBcbSa7KvYWMM8zl9DAZBL/zkdI+DLf+L/6ureL0VQ4rqL/2CYAhEyYkcxiom9q
+KM8gwmVvk7hwCFaBuIfDTA0IDCVRhHF98fh/NlPk5PsWsmj9sEWs7huTCJB5xsxLhgVRn7OFYj0
Npci8zAoQZ1Zvlnv5nHuVGkzhr6WQZ3XEKmjf11wQaUh+SDz/heR8enAJ8/DQneftUgJu8wqywDh
dxsD50UMiPDGgwW+SVMr7kz8jsnx67hw7tmAsMhxMogDqpjp/5RURdPVfoY5eqrtuvqqycIIJV/c
kA9y1vE1gFlSVzC5yhgJxTabi9t3c4CIOuLfROc9Bx8uafAw6rkF7OcUDkHzAwx/+U8AJY7FcAWg
noCCvqnofvIOfbXEAN4arLy7p7YzCEnoy+1VEl3YlBvFbnOxQqBgPdQBgO9ukcgVyNRRYklG3L0w
f9wk3g8ZEgHhJ/3/hwYIqAPo6hpfQe8hVS+OiIqGVvcQ1XM781jVPBIMA6j9qUTl8G7MDBQZ1UZE
aGslaWB7kJfYqzSFJbR+p/aOu6iMaRaGLoQ3EYXVk0AbQpz7clQ+10dDE1CGPFyiUUdUatpMV2rs
m9pKRFwlzwJKFT0wLJ1rl0IdLGGZozOcltXeOLTL8Oaou/qLpfChghRP6owFvgc7zbioBwtxAh4U
hSB3vsfyw0im901Gs0DyE3rpbpD3StKivIg6HnHMKWneIOlSjx9qp4tk29gruWEQHYmFZitcYa2S
BH8Mdj8l6+UCbYkSpYBMCUqEzADa+euY9PPV3mrkUqy8Z6JneOXER/lLLJuG6d4cj/gsPhjsomjI
WMRNOpyiyHqCM2AHiL9IhGnO/zRt8x6pxyZSC8+6oCMUVbLX4qh8bx98DUDQEJeugo3ux5TcYIIc
iyu9EqQIRGM4s+JNOMlQ/tw78iMkt50v4YNZeAC1VM1/6mwgPFRuEmGAxLchHeWkYhc2uauEU8n0
bM7x3OyE41R5JlTAhWwaVmDgovobWvegQY9uRdMDs508V7ETpY0wF+P+ffoZ4mtivkxr+ikmfbM3
bN+wJyylEDmi4mEq6SQuiiDGE3OAinaKTYa2GBqAiMZstWCsyZnbmRNTxxJ0QAw16j66kUUhSxCb
MH3bB13HziLaKxRV6tpXp2HoMaOYjTUxOcttfAforUlHohgmBoT1MFERVo5B9x5Ttc4UZQeQUDTh
oAOfwUrT00yb5Xq3PnivEBY85ydUWeNxUR+IrKRbQdm/tsvbg17/SLJYYAgK4be2pBjPtdqXYfWb
vq8q/iOlw9jHxZ+pGergcas81RgzJVq1ggymL6HQzUiZRiy2ojasWlCdnByYlsyXPAIaXIcCQy6Z
3fnGGutMdJA0iH5XE3GPZxG8/KECOqMGlEytamVi82nxoHjvAZZNRY8h436c/1yVo9gp30hzpY6y
Dm0f9C6c9lbnWlj7fsgisGrOR2fIW3v+JCzNdC3T94Llo6vigx1Ma8bsnHgc4sqItjRzEZpOJ8Hv
BKUObRIoREqM2h483F/zvnJYOZQ5vvUsjmKpfv6ymkMi6af+LTtPEtHyM+OT7P9t21lbpO/0AgnS
y+U88yb/bBBI7DelAqsHIdT3exBo9OsjHq4WuK191xr2oJUcCL8e/TVkqhm02+o0ys357YPYuboD
DXzlcMCvQciBvAiCXFSKPhSexc6wMsN7DXjFNr62N1PmjOdf5+XPWKKK3eYfgqLoaCA7ukNiu6q6
1pN9iOq4HX0eRZkdupcULwncyUehs8CYc+kic0sVKKrP/bs81DqJqIxQmi2v7CqzxVVO3o+dsmdQ
E27kg0Sf9mmNkYES1OlB8HiDp7uF2eeyK8dx6SEiEIpiVJhj1fsmZ52eOUPkMkw7Czmu6/e6vghn
MHg9IbgR8Gj20BTKhow4EJC2iTDectHSOF8oFBqaFyI6vGMkUNhoGVYxKmERh+ROxOCUgzrEzbsC
3+ejk/NwOHbB0vNgPv3BKVq613zOnOV//qIPS21btjWXkMypg7eB7Daa6saxcy8pfXWSvbmUxprW
4+PvoN/s3jGOXTMYp/E4luxvfjOrJpy+jUnjjhWqRfe2pIWATrwAdyhe6lqUQqCSTtz29K29zG0F
prS8nojctbvVCKGYe+NVh2mGBKqKIvecB6zGE7QLWkw4aQv4VuQJEwA9jCthHXcRj0vSmgKF7dHo
h9jzSE3a03vssk5/jzEoc8CMB1+Ddu6blRc9MGwGABDHdtFxFKkU4ea+D/MipBjplllObe9mrKvK
aWAI/ewcvP2Ksxp+Z5o10Pv2JSWO5+BOT1N1RZQporB82xXvC6o8didajVkDkzvZlHaYp2R6rAmR
ygxJxd9mUgXLCrxnpgLJekHVNYiEpvBi2kXvMFyhlhs3ojZGw0XGExvD9FIIZRqTl+XuHMD/V5wK
EKo4v0s+bo8GgNQsd0jpNGdoWmBwmQ1UBL5dN0u7cncn++PmwXqYO0SJm/9LYheInS1xEC8h6Ras
wssTs7E+7iDe+wM3FywmRTT5oEWW3OgHYj0/Dn2K6ne4sOuQ30qliwWyx+YqrtKDfrQ7ScQTynjO
Rm0Icp1mhVnJ91ET+ZX0MEr2xfPq7SFx524YgWmNHnWaNqd+Ls7dmNWQmSQVxUpfz4rAqcgDTFyl
lhTzoYBUKLgEKcQldyjOP62XsXOR9Xj+FiGWqZlZzNK718rrvVeW7It20cWXfmf2f69GzmlAT8hS
lwAfg+QwJgIOx0EobG5n9wpGGy4BcEE1QqyKdfq/Pov+kfrUWAKoQxH95JbxarmMcHeyzoZl74by
R0gxJ7DofjgqtCtX8Po2teUeLmSZYw38rmSbbTt/vDfj3Cfq0YXw4ZFHVfjZDguI1HL97Yvg7QN4
EwVoCLiBbi4RjbSgPjtp899oKqEFpYqnqGBla8uMTezPx4WPBzfwxDg+Jgi61lMEpQye7c8xPJno
tKCsxmg6sdMuwJnizLm7OWvKr6QdPVRV4haPYWNjn+htj4cve4PIJn4XzmxX9a7nWaHMkoOIDpXz
6YTlRO2lrOUf9XHiJBkk0FhkTCG4z1QjP9BikdoSBpGavkQhBpXPm7mqHQOr7vnbwUsKNrKrPoIB
AGMn/dA4WHXNVAhdzFXDpMgkL3ZAzIvlUcYLbrWUfd18W4YlLYzTrk6stpK05KPmqUMoya0hiNGq
3mhFg1tgKiohcYpfxzHiKWNiaQHG7k9wMzD2rqdkU1lsH4jpHykxMX9VDYr/BhRm6aM6aDHEba8U
Ya20rTRvq3AUYgJqYyuid2uqq2U/6Dr73NfsAlcwxGpZWVXEebXeMh64Y/u0H7xHbwXH0uRGthCw
TSEhHRVaXYE2XV7hhXfcwFCDizMLRubGa9mXGDNzhuRmcdunlIDnAXVbuXZnPrpfAvtsGdfx+n0J
N6z64zG4SxNgHZDhejweRVM+JLGNxJ6exU109xnC1KKxLKRdNsoQb+9WpRod7taCkp2j4sHwMve7
WiOU7JaXbQn8HDEDyLXfgET1ISV9Lc4//AvksZibPg+nPq7Hw9AgIGsKK0sZaKP+p+t7rHpR1uRx
8Cc2KqED+YnqKHygmBaZcrlAWshnXX/RxWqKrM5IKyUOZuOt9rhfdNcfdceHAH023Vyex1QPWCoB
dKPxd9dG4hYO8MNBDuAlB9llnnVNfqukGbL5vL9rnQzh8MXaqMnN5VusNBm8omijNxKYKczhkkKu
nFbErL+066sfpovPwtj7cIvJ2FaSqicZpBvAoQtL4wb6OV8mSLA/9VBim4WVBNUVcE8c1ot5qByj
GhdDbXl9JuIpLHKycgHphBgR0l3jrDekSq3JdoPeMA/4OF3aetipl2VVzXun4ZlKC08t4QXadrfQ
KVQr3lNTwXRRzBP9EP+jcdFoXo+EhkColg5sH0gvOFEa6MoM7PRkK2d6AUdBqxso6aLrUnay+4Rn
uzEXxK1zIr5tcgl5LsNKS2s1FZtJkYWiA+66V1cbLMITrBigjT4YXaYrBHuMon7eU3HStV8TBuSS
xMMZSt9k6itCuTTVzbdei+x4U1rPtMp4L3Xv/nz8ffbbpBB3ckBrSjjJQXp06llHJCzrkCCQDDin
xZWtk2wk0m1CWMeA8WpaYJNMzV2wQB9SZNwVR4j8yT94sMNSpxHwdseXajAtTc0CXqHAhf+qrZmK
ZdngnQX1x8M8j+fJ032iAEFY8KeZg7iUyJaDtKDri5c1o8mB++y/UeoAEOe5u3+ELFyuz2bqHQj7
aiKhkhfT5JRq/UJr8ZxrnJz4KY4Dew0SEIYvDA3UTbCH9ihxgwRKdbikdRTLbRu7hFu5GpsPB12p
a9rLp+0YJilubv0UTh0BZdeNClksjOTso9FdAg15jwG9Y+ZcrLiAJKzzHwVOoHMUEgVgWRsLvdtL
eH3qrVlBfq0B2Kb2VyeyiJSR4gk7viYj4MTMznI/xDw0nDmBnEkHRrYJW1YEVSY11RpWGw4+fUQ3
X/qjdPAreNkKDHRvR0fZwDpUW3DsfD/rzohPy5IEirmLtUemlSiQlv/jA+0OG4UuzEvtI0aw6Egd
wvTA9BtD4VKIRY+Wl4sE/x3f/Gzoqw6aIXLmbJbpkx3lFS9st0/1WVbPFtdI+A2+5hfaYIjR/eTh
TY39Gkaq6i18VaGM7B1BN/Nezm5DQY+Sr9CpXIgQdpbpQSwLg+XARNepI2027NdCqGN7AnYP9oX7
w4lkXf630FzmjDR8I3cVjsU1sP5WNbeU99AuW2Xb/F6FdDuG8/WNTgga0gzXt/j80upNVcGCKf79
F4XqO8NmpxBzgA5xmSxeu2Fkrv6DHN7JOne2cj5/6SV1evbIbezdZgBjw91eCRB6i/nQUitQXo3R
gz0zjRm/+JznsXVz0NmdK/VqI6lr3V7iJQc8nDQ1QIU8f5AdbC6UT+W6kNa8QW+hSsrdOgIsbfGr
0ru3C1tmEBxscC/fUIDGXeD/YMyaX1bphvGOXiKlmn+U/WX581shpAwHtc+iRFnB6xSmFEyvaqbo
WMeiCZb7Jq0Gm+8ykM7Zix1o7ctQI9TbGEGVuTKZWusJIfT8oz9kJzMjWNez4iNLFWKtte+XZZbd
pTH87MZIcPJHJMov5B89NHaA5U4Vz8Bs5Bndkzw42QGFTM4CgtFhvQflL02Aipm7FWe+o+s+Jo3b
Vc4UYcRfLAGTfS2Z6CZPZSTZBXpnZ1fTCWuLbpt1fskxlZRl+QIk/zCNF/kOVw006Xp2g9mrhimR
QnBxE16yNAFuw8FI1ezCYW4JJC/1VFGn+nucSKIf+s3Hm9aw4bz6DDwED+093SxGBm3kdPFWKgk+
Zut2SN34fYwx/qkcyJVDDFigsLTVY4juV+4nIh9K1Z8qyKIZVW/X13DjqIn1wIkb5CsR/852zZgz
ZWreTUpn7rRfrzes+UDipMEE/T6PL6QFh7bm2Z3OvEFD7F2WXnUHInxJAk9YGL00sz2MBhbHtlj0
DFdaWzNYL5ju21eeTRjR58t5QBXJ6hRG6mcwHiM/FcszQrPIhO2NeffS6bNkRUIWg5MUtGMxjp32
LZF53bTGWtK/sr7IiCzq93fjSSxqYHycEJJDMdyUIUcquNVk4FjuWiS4Y3ucUWimBysHc+87icHX
+ap1tp/yKLNqIvEvvnBzbQlch2zyfP4+LDgNeoC3qIB02avVtlQbY2kx/IiwOpE9YLNQUWkRabev
P3o7pnNjfwMA/9a6+25ZqQ/4tJ3Iq1riUM2iXqBDVQ2fbFm/jhPCbF9OQq1B4R+65CgZ6R0YG2Bg
IRGXCT/Zx9z+1yUTxrEAen+T8waCNBWHk6K4ZLfT7COtLhnOKx+baMkgXcdI06rh8fpXwLEw3T3/
lmr7FotCioNfTFl1m9YDOcgq+NOtoAAFKd5GFAnLtjJYxM3EumI0cHcj0hCyEw8uGKMorZyhLHKl
JY3tXgmcEVenIfPumtBFVVXHAZ8rReONeotpUlrtH5L3Oeh1+Ob0S+RO0tjPjkkiSnR9QZzw7Ban
M3RG4EwWAz3LKjK0DAa8eUmbw9XCoJG+lzMt2aTi8t+USJfjMnQfdXaEV85NZVi1TsroTzxarO08
wRrsoHDxgq7y9qAdzRZwEe7z5WSFbYKdfn02X1tYLgDscdXtZ0PQdY6aZuZ3ARYatfUny0BcFGen
ENvn1/Ty5j4o+/eMrVilDpbHr+yjkk2DwGzrOfzzJ7FVVXXRZx5VIjGtffKINj7Dk2Kb4cqOw4IQ
e5i2Ff+W+xLslifeCO6WrvKiEsIYavO4ulG1cqd2F/8hXblYGBUlaXj9P+ZvsADtGrPnoufFCxe6
tIlm/ftTgHA1d7+B2yXvZ/DJdDe1huUUXTtQA5MjIeDs9jGxbj6HN56RMy4ZUkzerfaorOguwQ7W
ylYwj7iYeJQJILGrjSOAFv4aQWz0EovzPKobZweM/rMsQXbf8Gi8dcIttwnvya1JdEuuq+iIXdfs
yQ3EOsBDi2rPTZi91wVgFLjJXeeBcMSqYKAcKPyiV0btN22FjOdZhE8ljUKd9S0qZYSOlpYSMmCA
xkTSTSwCj4xsaV7teLJM5qSr8Q+04wEb79agRz/KTsvALPPL7xCsg4Beev/32L/RxN/r37JRY6Kt
U31hv1i/MakPLFFmeHjWMu6F3YRMDVcmV7t6IPJ8DARFuPTjBvwEoKUBKOLjIvFlR7qFZpzGPPXR
QwgRfMXvjDsAwGCekKegfDaKVC4k/xjcxWDA2AbSg4O+a4sp++DqT+ASjJh+WWEKry8Lf7BYOh6M
A9P9ttu2sK+Q/4bWrMxuHXLQsUTrOPqi5srSdiws1oLUoirxnQ86JQX7lgpFkr8YCBz2laCh+hJf
ktnRkBmrozHzbx1F8GHRqO+ptq2VSImg4YNhqwT6Qjst1Q9PnYXGsNb8uPEBL3C7F4CRS/5rJ+WU
MdtW1McY+Y+uBfzLfeNORRJ52JuPh2PtTygbaTmyS7+R3EFr2X6mQkMLdt9ytaWwjDIAq1H8NSw5
CMYmvfKkcbq8ptP3qnAX7EOx/oksgLsI3ChzA2vMC6DHF1S7OXFL6gtOTNqG4OZF00n6iyUG3L+m
YkIqLSvlTVibTmg3PQt0yrh97nhgLkFm1xuCnYhN5RDTw69FYLdOqpC258WutxFZfVYnFcNJ4J9z
C8zuYzBurNTI7L+OZfwpbgpsLR8SrRrcOrzNsCD5+eAkfiyPxDxvKpbDg7/iycn8KvpOLrKxbhya
E5Vw23/ABuBW6x3cxi6ic0SNl4+RO5KcRFKZTz292jyoxcKC1jUO4gCxxwztRN5NzZo6Oc8MU+F+
KGMMAZwsw0fdjmMOcr80GUVYqjDXtsJSs/0x5i1PdSbpXCN0tXun2PT4HwS59GLNplABylrUp/o6
mapZ+3xrVbJTIwUu645d8hfV6aDHXFywIQUNHBlPeJkPYGU50T1eNa49npakO8TzqTSPmmm8DoCR
L1GXb8H0CUtKj0fWP9AKnzMuXFyJ/ID7RdWAkjfohXUmSOaTzbguSdc/LzJcgtRV5qEDr6C/31/t
2st3GvDDPcAvoM5YdkXK3u0SaQ2YXHnD/hby8SwxfUTnrxah96DlZkFJd6raR00Nr57grVC0a1Yf
7kbvMxMzaHxAJz8Ku3vR2U8aCt3oxP99LFBAWMocQJF0SGF45MJOasw6hsgGXZtk1Kh4epMhxgz5
Q3av56aQaDGNLWs8qvUaAnB/upXCsY/X4/AYF25a2CxRr8curumpwJQ7k5pdVXhtxc2Afq0KKa1N
xbIRTuYhRpGu9yzR4YQPO6t8StF3DzPKJYgs3drp/PKo/yQJDj5JS4V9OBaU0weuwPLtbfCHM/4U
k8c/L1S787tr7wXIHy34p9/ZTcHljkmigiNuIdt6agx9fqNvp+Fed4CcR0gR/Pvtf9KFy2hey/P7
YG3H/mlG5DC2kmzkcdDjjKdMy69ofyzydhfut8TREk3lB6XKq3FaT2oD6fSK+tjRgORoow+nP9F2
kPUXxukRljUJCiZySkGHji/uXUwKBZ2HDAjEw3u5OscYEwdEtkvIo0/SBu2FwcK7lGPsMAtifuug
I5Z64/dpKlGOJ2YMf4nU3sFRH99mUFN4WwFe6OfmruSdo6PkiAdUwG7ZbRvUCHKHvqF+M9+FrS4N
14oc//0E+y/MXw4KJ6OAHavhRHQPVuSqUgEPNrHE0olx4gBGX8f+ZnauOThGlpGGkaPAk8lMKeeK
iVYMRSEkydDSVHyIggoZaf9HT/JnDgE9ZOql6BAAQ6KM408EWnkwtemvcKXhHBi3JX4XbkiOWdv/
HLleGTinVAfi6HOhumkpOBf4m33idg8Ky8rPt+oeJ4n3n8ut8qaFBou5tBUL9zmUYuRHw4+3pc8e
LoKe9z/JZ9bWkuwZa8eZaYvSUJodnrvCWr4ya5+33HpAJU1BwwsBMll+vzDk0dnDa1zznIUCjbUw
ec6Dc3MPiQgnuG5WWVzzvHRds162aB7xhh5azfonek5fSP6n0Z4aznxL45Sv76z/NXdSrq2fk/Bs
7WA7YK2IQRmyBFqdMlBYS/3RUHElOR3fyn7/VqmCz/+NDWwTxqxd+/cY5BLmVYwdYGm+PQr7deJt
cpgxIy8PpSb+et0Ref5maia9rmqWvqY6MIKDx5Mbcs6ruwmkVgKaAZZsdgdAAph9xNf3B8WnjXFq
qETFQJVAZRGJyJOFZvt3BX0saIXG15t9q4DaJQrtcVH2OfwoprUcy4N6M4qUGYmf6Rvs5ey6cHT2
qQXGWj6HnVGXA2/JdWdHe5Jv4sbaG3VnqW+wv7AeBTG2vz9xx872OsdHWOjuwHxNL50Rj47dhv6a
ua7cd/aFlpxyku9HyZ0+zzFfeU2VdGt1vmODGAzLtTD3bG3vzy1kqXZw6BZQBYYRWF0T2RFUgCq9
cpj1NukFZNszalVM4Wx0U4pi1zUrYbTnCBXQaYRHxYZNQI/VKSTXsJswXgqx6rj3W4/vjIQW/9fD
bAXqPz+448JiJTzIrFMyFJouDm+3sVPh3vWuLWVy1uKLgzcdtIAOd8Fyj9Bmj7DkrzLwvudXD5SD
vSraEm0F5W4t02+AMOpIR04f/Q5331f9YsBnKmBVKftLa6tZeDcgtYyJNldhfbJj6teTBTb5zWSI
bqZJWefNj1UGct3Y77lzn3UFmq7GgKKLdedtDhCgIrxIvp0K2CsDoEvU1VYrXcIbvtsbzRI3fvuW
MfEdLsJMHrvZ4FNLe/nSSNC7N4ffOgFlIwl6+M4y7WV55a8CtasKIOK7J0/yYbRgqvdmaJCFn0t9
1OPgV8kkZVnm0Qnt2Cm6YXgNGlnz1/Xvn1z6JIh8HExnmJIFOJBUkVYrfRxwbBpxvwxBoV6IAVbt
HxM7BhCJqmLi5p9+AqCh09Ya929lrtofmLfUr4heRFmeCPA1NRAgPK0one8x2i3Zf0rG4ogrnHmA
Cy+2IdHN5KHaZSo9b8HfKQy/ZiTPmloZBoH0uZXhD5izJx8C9z8fjv6aOZCf3Shic0KZCO7A3PcS
t2Dsh2pFsokbRZJjXevte7zWd2tL9zMhCDRA0XRaAMDzb2qzWtxEhA6ACQ09iG51tiqfmccpQRJ3
3dps4E8Zh0NM7CcknLFrnqj6WBjzKalKTWvxRtf5H04NkhvjpcVxsgbNyuv2Q91ZQRNnsguYK4qv
6nyJotEvzGq/NQTYTqJJEn6r1JanIh1cBK4ESZL8XdsKavUzCgzZDOMOSixgBZrZuTkWEH1NbKuO
KEnbB3g5UyehsCAkdMMSQ6KIJcKd+y07TfvnvVVqXRb1jVYjtOrN3KbVk0F6xww4EMy0tTemhR8i
/XUlurWum1clKgnap/mCpQGGy3+SVBupl74oAhqiY9AxA/9+Ewf/Oswj612h00Av/AtMbSO1sCfy
201ndzZiYzt91EKQnGyB/ovAxNznDXsFjAMyK/tIKkyad9oFiCo6555MvHl83vz0pzqaFs5RSXQR
eeQ4cg2RigcHmuFD08SgQGw5obPScinhdRvuxIE3Ka3kNlfrEytgdf9+rDTTiWg0OgbJwiLJKpYw
anGOmktR0q/3thCd56PiUlBQDHRjDWUIFTbGva3vJN4phrbnlnCsde+GLdDm61d4HPSeYgrZYMpG
To4fwFV9pOjxI0xY1Ie3Q7FNOUUcghMCX/P27hwQpb9S5dUeZDVeoHwxq1k9PEuRMAUlmyifB89P
OXvuFFfkLSs7Cje2MnGe97oxakOTdK7rr3wMFhvLxOjez+sm6CnswupS6nbYynge0FpeQys2SCeJ
0FK0rMoIubK9o4wr1HZzn54rBP8/4C1wA6AvaDmvrG5EHj8oRp1PXJoyW2yK7004xWEyslvf5EYf
in2c/K8aPdNUP4+8evc6UYCkiPKV6IpswY+41D1tRBButrwlxit2o9EVwQLtmwdNLJmMe+MdNXh2
tyMWmAqKP6m00QQ/84LbShCBs++6UEs9ngQH7JPa6+DIHZxmZUZjWA4KJNaLOIc+8XnWS4XL+ELO
MCSNDBLtmgf76612YLyCD3iZM9N7vstLNasPkHrpftR75+C15ysDhPDfHdcHJk0l/+cBshxqNGmX
qM309GRg6NuAgBTrAV8ZECLecu5yJSQi1R4Mv3674tyEU5ZYPUZhvETGdBxMuTwtYUKjLKzrpfK1
HSUHmm4LECGBjpyUyHKbPoETcymo19YJq2dnGztJpnRhkE1zPd0PGd68yVnRURfy60zVWpTSfpb5
B+9V99VzG2dtYU6W6ZDWKwT9T+eivSI1ccvixdv+gLY90Oj5gixh/mz11xmd73AVkc4MbMQ7E2DZ
i9Y9lIDJbtHA+PU2x7+VZu4CQIYVZOCz6KsypCX6u2L7Cs7hw4v3kFa1mP89k0sj9pu57kn0JGZF
JamRTc6jSFSd5jHNMWgduesKSwghYGzeWYSNHrx1RDZbHhfxemoKvJUs4DdxHQpbmSo8T8Hrf3gr
w49faIQrkHZOkeelmHXTceXvUeINDQ2oVgZkZxvuqbsHcWy1a23UhRyoDPk17Fosb77SDLO93Nvv
6O6I7pCxxY/+d1CtmAzEqwgxoO2MF9qXIchfyTUdD5CBmZLeGrE4+CaZLXIi0uAeHg0kmSsuZD0M
O9jsy/noMdi0MXaLBioTK9cG8XPeYhA7HihVsvSwMlCwDrxFiDq5ajaJj2ygJC+4Lyx3H51SWAYd
Es6FL+OYBQSR7wZFrbm9DQ8vihLmPny6IxLXOVDe/qcirWhWGCkkMmBmr+CfbnwEJ9iMDkIAaW+G
RK6p0Y/xFaXQoPlPRZKn5RgCWBJvemGPRcQ/phMgwyxFdSf+AjYqRtEytXVfdStKmAPdUdys4JBj
ROGhzSoSg2ZaER55/y4guzeECtP0MNT7wWCYhn+i7gV+z9Gl0yn9BAFCxlC9qhFz3mDC51N5N6ux
i8dh6gDQoxb9COHB5iWH7NUIpHVBDzIkz3j99h8Ddx5ZPVnFPtc4xN7lZC66SAu5H+UHeSJqE9/n
cL8L8tVbRodEHFCc99IPRlQKW7BFmDpnNeTi0wTPx2jIQTyF+ryZ5vNtUg596aOKYtkhOXRmxl/8
dCvXjS29puVThAefamGgY1xCryPZe7HOTeP+Zlf4HxQ6cZ5ndnUfAC7shXzMq4Oiq61vlkSR345E
gb87h75IIOg/jwSpzngXyKXhc1beS5IZ5McJ+PIHKhDqRi/fSrs1F0CDPGSgFsfCeE4W6RPjJ9Cd
kmr77xflGmICpQAh1o2LWWw4XICxWeewf/mMKFbjyPV1KqCdnbrkTSmjuKl28xaSqaG7QX422xtP
moUOXkSgMnHwswW39Wra4d9/SeFXLXw7ikkeCxJUD2EEhpaCdcsOS/kYemHhOdhsxyZWPAXQzVbI
14CaczdHnVxCHps4vWm6OB9b0lUlKP7UBRGLzejMU2NPOJH2EgLQI2DA8dqas0LfVQ6tgeSdblQ0
3Y3FUmtW1MS3Mc0bOy/ZMlLjvfZb4N1tJq581eGNlBYwipG4bTfRNv7fcT2lQ3vDI5WXDDJRDvLZ
W9O/u1JNl6d+ryZGOUL2W/JPOJ3RL1yI/3FHIUPnx6nZ40A9+bIzzSaaAOJyfTz3miDqv07/fPBl
a2KVkbrhsgO7GSnZrHVP3uQiuBJOE2oz7eyrU5wkXedwHeVxFgrt58Hc8ImBM7fFeov9QrRRIP+o
UDn5aSrNIDaGaMfO/n6lOR8cg8RGFwi5sQj9ufuwtczueKR83WfA6i+ZuhrX6zpMaJK46NY3us5l
B/ElRNswjHCONw0j3tXw4/TiGViTtqmmRNqeh7k1Xky/c+MpzU1OgaoSs4iGlCTArXD4gt+LteST
H5dmYF/fkUiYc0Z+vcdMfrK9Cpb+kAAjVZ1IG1HXCCbsjVxivomEC2aq1MF0+P8wuYXCdlgmNlXm
8XyjTwfkKUEURJXBW4ELsujGznOd4v2lsF5M2Owktj3y9qAWqDtKY/XYEm7pA2BcHIxR1M9FDpWE
Ln3La5jQcFBxi16k00o5RvXuVEfDR7G7f+fKo2Apyk19+AFUcixkTBUdQ1qTMRsbyAl7BkDhCzxw
dMf1SRZWeDHC55WTLnH0VGwZMyWSm0JVMbZzjtIOLTpaOypLt1zbYlDOZ8ohoq7N8pEhV2tSt+le
cb6czNkfKsK+Va89jQcZ8HZlhG/KabwlerCFh1vJV8zEBeTIcNvd7zNeOwh6aARFytHq9iNZimZW
Hx8k4OTg40plBrxfX3JJB2VLIPZ85447/lJREfgmBqDROWQrAHvjlg3Lt6Uv/J/HRdWYQdLEL1Ei
tCgABY1rpAux8/ImwYfnp08xk01veWM2mYP42qiHorGii0bPxsbyHi5lpwP9H2/+2qSBl2br4hot
Ea1PZWhQIe0CjhQa3uH/o9KHUTV7XS/qDJjbugwxJcwPPE9oADt4bxRqnFIH8qTeY3MAYTuWU8Xd
Ev9WAw1lb6gyvw6vgUq64OF39AYpypfJYYaoMVhgHrurGDdb0fiswrsRXnE0Wrk4gpfuAkDQSZCe
zxtte31rHfXX/dTbUQ/rKo8AD22eRUcGsxiXV/yjOQRszc3Hti88d3gcfkSfjDPGtCjZItFQe7XM
DiAkJZBHLqGehCvO14Cq8LO4xz6qgvJeO/cJQjloReq6uu4SghcvHeMLm+gP6KajEX3+tzaDDgdM
GHgSRZKd2t3R//Sr9vc3ZOI+oIzpT57BQjpdPlOq0zf5fz+9ofRCHiixCxAe5hDqjqHskIWln2pe
VZLAGHB4uAJTVnR2B0h32RaCpAQJOdDDaBAf2zPOIitfQGA3IlJD43ylEYTwBOEVrjnFZqX1zmnG
Jx5RUzJ2h7t47lbhctz9y28RUNN/ulqUp0KfyROR7gdcIOJRjQw0oObRu1NKkbguRd1auUTKPcD7
OSm5t8oh4tFbizAWTGU2ccwiuv5RwdrCPwmatANJueAxOFniFh3Xnnu+zgaJD71rTf+tpj2FUtHr
iPIcDN3gFQwXsACeZG1ObA72hJ0+MCnmqDmT6sGcdvCQZyd2eBMGUL9Ayb674rq78GJBG5SrH3eh
yd6S7VtxXt/bWqTGCqPhjuizh27nhWbuqxKLzfSascokNDYG2nTZrEW5Txd3VhyV5O696y5KunBv
CeNjQL7zar40tpe3kZDj12CH0hwxxbaTWopglDGlbC9fFFZQ6QHNl+JvpWi68eQ1UxMJZ/2WrIGj
u9G+2I+HkGVSRWjfmjJEEaIjTWK1/ojhciMg8NDm3Ap2C/xSJbJOI4fQ7S80aleKNyv8aXVAJM8V
Gf2VJyTTp3DqwFO2agjDFOIKV85K7jHsF9kvov77J5MbG7INyEE9Zgebdvg7OEdnBq+ajnYI6QlV
nymNXQbSl+y+e2tkDNPnBNyMNBv+JDnJ0v/r3XPx+ec+lo72kJgkPuewssW0hMdWU6Cm4bjmY6G7
IikDy7RlvNBAR2pDGcmgjFS73ZHvTHO+HdOJ3hae+mD8bh56m7gssEKfstI3Fp6RFQC4BCbGepTD
bMtcvdgm2VY13iCYiWOC4rVXVvg1Vf5ex+jlw1UBgtFAdr3ENtL5QGUK6WwpI+laYYwUWPTKZevw
V23XP0NHwmv8fGxw1c44k8+n2tBCw8ozg8gztbfldJzh/+CDAn8L/p9EYQ6/RHCyhWR1J7RFzErL
fdwzdKUFve2PEiuGibg3YtTMITpb2L8+g/C0/i3z+ExEX7tAr/oKdqVAQSt3O/V6ihPQ6pJypjjl
kVhXttDDqYJrJ3TLqouhlUjom6UQS0ht2E64oRtsswifhe/acBxrbJFOQz4I/L0jGBa9c/b9HMyK
qMKU7gBk79Qnhv1pFHj2LbqwmRLNetMt8AKXhR/8HmGmbIb+IGnv6wgl4aidZkRKorjrAvPNcXEq
qjGCpmggPTo6QisbRWAPlhe3Kebq8PTx9dzLbO6r5Uubi3EE3j/0BypX0zhU34XsEw2JNEKRjKJ6
8Wa7envfpsRWUFzHhxls8s730nFzFBRL27X84YEQpVz1FoksdKW2IjhocxaMfNS6b4fNgSIQj8Z/
53O31zskTViMQtDLFlip19YgGY0LPv0uo8i70j2oKhcvqUwYYlVVmxs2pJzS30f/F6KELhobA3rq
adwyY4ZsGwGsJsBbicILQPJs+oKRj4kA+9rgeDUAxCQVvdqAHacuCCHLpDdKfPjJL41Qv7aKDPAI
5WRUkysRKACgoGFkHizcv8Lgptoc0B1v9epcFrRHWI+D6wJO4qQFaS5hMvris6jgxjTADmLA7oo8
PKJujCd3iVn4dLqZzUDXz9M3Svpcc0qbf5749+pkSwIr3/AXBMEaix5sxyqRkF6T2wtlEBqqSMPr
tMPiZy8nGCFYRc/5TCpIc73TAbs+8BxvAGgpCremjoQ/u4Ghkqb2utUmh/QU5hovSMrOc8j1xo0a
ZAFj83Wcj29jsJ/ldG/jFiel10s9k3xOtGlpaaTRl5KG7zrtPxx6PUfriwoQjgIRLbFYKK9PqFXk
eQfCyX+juWSH/nF2oLEVCvUQhn2lBDHaE4Lg8EjXWL4t45h00+yiLFvpuN/Vug85Bj8JFaCYSCPQ
KXVGTLhR/JjM9HbvqdXI18rP+gJaN7toDHJtuKiAQMfB7NM6/UzTqbte/BY2ZQnm05EtGRCZv2dO
RsLFtZNc4DGfp2xSXFdqxlq++DZ3E2a/9LEDkwYIEPRFhxM0Q56b/N1gGJP51TeC1YAAcvaoxJAy
Totj5siq1fobuW8Y4DwL0SVctPdKTtOFxSP3SJX7XJFLGv9EcPg1sNPdl4foHQOEoNC7IiTX6ChT
SoMGx5rDBMyk7VRIqYvbQOfzC6xK73OaGNiD7/qoM/0SofS75h+YQVad2pYOsINpTRfgdzU23vbN
U4sDcu1VSbGomSW27YTSInutm1XpBa1fxp/ug3xPvbreu/8UH9pSo8Jb7HJc7NysK+VUYRMK+kLU
8BYMgX1Z5qSNczHRIM0zZuS7emW/HpZE+xm8Ll//btkZuqR3FZ2EXxgFib7liqYmrHcsgPv5oFbb
E/TvA+cjZzWreVtEWIeqaM5iMXHW18y8AXL606N6kp20sscUmW0g+A/ha7unwIGrJbzUAdBwrt2k
WK3A8IwTebfmKLC4AC2yNdfsiHgQ3Gwr0curlIB3P+NXE6nZyTHbto82CR3KRgJPETlBtNKQmiF0
CwgBMzF7uh9XHRQMKnraHcgAjNKALgHOSyUk/5m3fM6le5pEOnUgH7GhIe/dsc1btRZO55wVzGnQ
MkCHfJQ9b+zvpNqpZz1e5ErE1N82ZmefRwNx3J3e+zruZ4xVKhPVu9Uc/5q4iPf2Y1t5yMtTSPrM
UIzJmEQp65s8v1Qja03ypiMfN41mJnLyLB2IwYv1g0rRLEPMRZ2MjDp6c2T+OHrkve0yLfc4Js1f
x7Se7+EmZaXwBGRhsFGIPhRZc8UFIN5UgtHri9sw0PHCqD71ehqAcKlL4+OMjmNv7KjZEVV6n8rQ
fxFv87+2kS4yv94YWXW79Ks6fuSGkEXiQ/YuOH4GX4A3A5ruNG64evZSXtMcWIZ/liBFn3qYYx7M
DCMzC2K29V86FdfS1nIP5skjzaTSNYIzxgReGPhR6RY1mEm8vf1h0FI5LKbTANrAw05jbbe+TUjf
u3b5N/HrIeDg4teTYdKZC5PTo2kQgjg8aAmxRny0GACuAer/o8zeYiODtaM45tgBl+YRXUI5BwAv
TITdHwFp3GRQKgkXswWDr8f67VKgp4KcaMN2zAqVp7/SOrMZUnbHLCne9k0JWPSxQrQM5hyhuSqH
PW1m8qvZbKw2zXYXEZlzjVfssY3V35BS90GKnpDCiRmi25VPA8FmQmczMpL4AdyxExfAyoTlXc1i
nJRDtQhYFlJMZMnC/A9bHq9/fpBl0P/tdrBp6NY1PTZcdhKvQFMr5kl32krl8KmyxDAQIConGBNr
YxCBv6PYBUdhAQ6SHFqwdkD2ct68mfpsjtQ9KdA8KCv0QTGnJ71U4ONV+wNm8rO7dsHCPIpzP7hr
EFKMuY5gXvByGssqGBdfNfEAK6Ki3qFpmRg3WTzLqAT88WmJ3vvsPoNCIKMeU2uHpXE3VAgzj4Ws
Vq1s5Dd/FGO6ikiEg+DXij6PGzu+A34MbMfvnOft5T3g09OOXCjChOid5jt/t4nXYcqbUiKwJNdy
szDTYTEGpDKxRkmU9MxTeTiYkyQL94XtBdbm/SmYhbUYQVVnVJ1hOai1jXDVlxqZONhXPejtic1x
VDig3NG5KXnB0Y7H71DkTKmM853foAOWSCBFkADorpC40q3GlLNYLt9cA+quV+26jZa7AZRj7pUT
V6pO4VYyJ63ZLVVCk4BvPia8t3Jvgp8Or+su5aB5EcWz2Rso2e6ay3xl7sIjko4sq3FC02qTMIQq
XHpijKlW3SSUp0QRFtPvwpEupHWXojx+0vQHIGenlzsMfgf+sGdXZZ6mRfH6bCAaGgHTWKFArpBw
2SHJmdtPM6BLmKdPV2Juo/gdoSwdVHVYqu297pHpyC2evbAO4WwCicjCTFCx80iQQJk0HbPrv81/
bhYWVorhZdqkWPcVyav+E0ghp8fV9B8g413kjktsErc9h4XLVX9yCWlCbIFXANM/Pf3INszWe6sU
Aay311zENeZCpjtpLsBgkmL0d2WXnoZZ04DiLMalNUFeC0LoQKJxBYQe8MahsZLpGhmb9ZPFOK9T
H5rXbX3bmdbdInwZvSxbbPX4G+MZ74AZfQ8hdDli5HJfGbAKXZSjUFSJT/tYrfOF+yJyOQJGSCq+
/fd8fbbLbzlUJhBvB9GwtzRZTEyY7H9WoYaFdTxaHlivHCJreYTt7lfQniZZhmPpdThherGcimy0
Z3gDegW5t9PTgxyc3g1pnjK9B+Jz1I67NYidXCXfTGmlLyUoFJ07nVTj3yYcSSrhz1pPpJuN1EQe
ALsgfC2cA9xzqI3NngfuTLx0rlZElky4gtzPn6q4v1bd7jTa4xTGcMUEFf7i4Kj5kY8Opc5lY11i
Q7MhVfNlu8kEx585kYEtHnsB5q2irU75E8Gm+wpByMImXWUnaRcfe+gjmmU0lotSOvFjHmK9fkYf
b+MnWC8eWoylevp758/ghDe3fdXBG+A3O/K9QozuCJhfaShfxqMwNegDDS6+TBaNQhEF1p3DiMrH
ZOpI5MXZREC9N6+HDKbWGfmkDEKVB50F5btaEPvGGnWxHF5y0Ye48x1nTEIPWA6moAzATPkTy8dg
1yT4kCYkbONde4xJw2oJ5+OzCu85L7evhf1b8hkQPIIVqSm77zGio3ehM82ONeaUZfI1BIEXqoaA
h1loAVS6FUxjeiaJ2xQJT4JTYKrqSH46Q68t65TG6V5ThgazEyWQlXK++g4fYaDISG3pjlHu3pIo
JbfAJx1W6s2DAKOHvnJpUy31CEAm72/uj+gyz3Fky/kWm1r4KaJX5cVAKsFMQ4iJDA4BpdfbVqdx
5g1GfAyxvBMCaM4Mc0WcehWKcmTVt41BlfULIg+cYYC4nUOKf+fdSZ2fZgljo8cs+lqwgcKiDhiA
1Ngr2VaOhl0FypTUFx727g6+mnLn4GREgBc+M7PapPkrb/wneuk0YOvSME6/7VgADBTrFspnLbfL
kAxhA+IFxNAe7xOMwpAfwH6mfxpYbj8zeIffOVKJ+2XhkzU9m9sCF/7hiV1GE3aTk/WQcKwvaDnD
DYaQFtvIbQ2YHbzjE9bVy1sqDhku+vthw7i4yWmPOp2yaTfiBxSaSHIMCJGNZi/W2nS9LhPp3OFM
CZcxcSidrTCP0o8MV9NTk5SRDrIGdRT7Fus7n08OdX8ApcQL+jUfXNGIFCM4RMs/eBgIIte1g0cK
JIMmuf3LdUnjcPlgxIWPqtswzN/m7VgWclXQ1u3gYhk5H7w+MmQxtk+zRU4uvy4SDK9/8hjSaF/k
JPZhJGsfuxuBQSmXTCbMX5IXdgm2xudK122djWgc4CerUTsCNhtfaV1gHdT6pJtCtlAk5SlPOOSQ
d2ZQXo9xzvnNe3AfNvm/s85mhPTmknc9Pfl6xUJne+rpJeBJ5oLMGb5IA0NxZw3DkS1eha/PplM5
SnV9TLeghhvkqc7hjw63reDnWPQJoDTG+V/jXGj7H+c+T+EVY6id7RJTXlu8a/N27GtGHb6LYZZN
luh7rXmK7isMGuxtpTtfiZUj3wM3vkC+gWZNIRino264yVIpvAov6nmlzLF7qry2oK238vJYuD3Y
0UFKjSSJnhzlFgnDpgnpGzKYlYPwTyI5YxE/Sk4Vzcbave7U4y39s0eaYjkgKJLE8+hSsysbTAyS
fM1ML93MEmMbnWupeeHgwynzmeDDTEyxoGZFFrraZYrES4ym2a+7verU9+y2UjYYaKvaDQVNVmkY
DVwv++dBpCtYHT237b7122q92CjE/KbIEqn+Ndh2CxwP9Ib9XmpBRRLMwFykDu+bwSBwLVew9b7Y
JxcDL+bm3eEAqh6EgjHN1do2zRt5HsK/pJ+HWdigziqDPqGlM+I+Pw+chTNId+zOK46Gobtodh5+
sKiJy+VRVxifMoW7/vZJbk72ul8YYO8gUQk7jNboDeBpTjn6iW6yuHwvw32na5F8K7FTgpzUkMXl
uteC7mFHeUJXhRqbT+em3o0nGa9uI8CBVqnukpziTNbRDN9yxuMivG5UlNl4IeT+QjU6IIjOcCjv
1sQ7EQf/lfCLcrNqnBQ3zEncSor+YDQDejtuFISrf36iHDsmM376/wcIJ1LOfvIr3KMs3SVBvkjq
iP7ixYNQmvEfuJyC7dd2KMrVDCX5/R5M2LXY+GGLDpvWtj0WHgPfkJ+rq16uZNCfDPlmceMBo5ve
IeGGBn/mmPLUWwugosuzqY4x1A6hccAqYjdi2TVa+EMxf/Sm2RF2288F++ciKhvwYaCQHK1K/UGv
FN+ZeFzQmB0hLf8A1Mv6AI+uG+Yti43/sp60Rrr87Yqxg8k0dZUnbd179+Erkl7o0paOmPFyZ7GE
B4AE0KS2w7AGlmcHmmk9qqN3CYT9eTXqhBUW/+4TiewQFvSyGasYcR9QjkjELQe/E/fJ5YxORkyw
gLnaS2FDX9drNE5+UpxvbAHoreG0t9aS8etE1Ka8VuwAB9Gf6YPVJ0YcipvqsFrFi4w6qEY9Xudp
d4+fr+SZTFWjMW1XpMRNlrSS1W3y0uEAFlgqt7B+ufLQprxyp1ltvCEK3apLN+sMaALU1ssIK9dM
j9/26cDg++ewHxQD/XzHMyReL/6natW11/RbAI9/GAmIUoFadjig0LiAYYRO1eoxSa/IwtOUClfB
x2bEf95WHOtag6p+r0HkZPD/Vudd+k0tL1rHmta3GmbXhPnfqf1tN2gV19j3o0AsmiXC77dEJv7d
1Ml+HXAOctFn/tekmqtI4sFP5IOl+nEzD2KTa8v75x9scuToVMBWiYCg5OKeXhN15j6U0c36J0y7
YqeY2UjRWmGA3ZrpHjnLQNWvmQkDmzfcWRBSqToohmUZTJKEKd7m2rz1pOZei16AWsFOYGoh80M8
yFsTCZIivWeMj0l+/LjIhWaeM2Pm/M50anzzXWWPuZiLajQF8I1eGQYaEHwHlC6aP/vcWZlX4t2g
ntCzbaAEUAX8XSgMwNGENIT2pdRC8dpikcEpPlZffKW2VPC9unput1SnZVfUoqOsthqC9fPzjEt0
wXdSJHyCdEyyMl7AfMnVZhGFS6LQDpJfbtKMOLiFZfqTPZ4mQd5LpVL8u0M7HX5exJlfyuYpAlK5
pVSmji9ZiKke3QxIk6Z/Y3fWVi5sdgSMOnZy4UPSXH8HJ5H7MEH21XiRHN/kqBslkDLwH3faAYz2
LJONFi0dgpK0gfPTMwhmLlPUCYNwN9FrinNza/Kse19JA5eMilrwOFNa+Gvjcjmj+Q725x2qf65+
4bPWxMGckKvj3RN97sjmV0Zx3+S2ZJJFXBFPd0mFT8/+3B1yUyJbfy9MB9MPj+CoVQ5725Ki2xuz
+5LPlYCab/V/aTXrtWnEEvbakvRLkYtGUtr4C0pU8vJHc52zvElUTV3zzYGpQrjnTj6LmZ/3/vZC
z96cxWGIT5GNYjtK0IeyDYOpBYFJUhzw6rTPiPiygiG+FVdYRUdHhhdeI+eKiBGV5ulDwsYniP2+
/00pqX6QBJIWrNakqCvw1IsHzbYoJOnzDHtajFhv9l6td1QRTMvSF08xfJ9vOMsoYnojUuwvXqAh
2tN4kqcF83I6eUHtgVGjRDDr2+FVSQ5kIxIjlcm+avV4hb7BLz5NK6MAWRqGfDnb0vDvRkr5y1CU
GRBqKFj7SQCzkZtBBuxc4oQ8VU6TucveCFakSbie+x6nPfxOwMMrmUAWa4cV8EvcEBIizwVYSe2g
tZ9hb5mWJ5jWdOuw+WQdkKaqrCyl7Pm1XxLiDJ6UIEsR10H46O4mgANrIaY1nVakLqYmsJUgm9wD
ZEUkd9Y4VvC8MEVor0g6qWPESIITI7YyfacEI/Iq+bJSFx2ccwBfH8Yerj1aa24Ov9i0rcery969
Bjl90mOXw1R9LZjpT4eWthfsjKTfgAKbu+/mms4QfjdhJRnNCzhBVeDYTahwnjBMAIWe1IXQgHat
pDtvVHShHqf4m4nwdZFLrAAmYuqRVmnv82Jtn8Qlz57Sr98YHnvTulovO4WStWVQnlDGNnlOuuhm
cv607Ni0OmTYN6G7wCdkw1iUp/9+XWrnWjAmMbIJj6Epq5ja01Nz07le5RCZbHTsZAhCm7dou1Pu
iUV0HMIFbxeGeeyNOJXH6F+PCfTjY+yTRTZKkaDgX0KG+E0Y0F1ahG6ZP0DsgOFSTp6xCgCx8Opx
PfpQXywHVBzV6Njq7kyIJhQKHhqu5QQiBCyqKcNVPxaIJDDw7I3jgTaP5UtnQG4NYkosTSnV/cwN
OIIZA5G2bOgicOxSCxZ8iKyHrulMGAGcWuZpGnJn9zgFhxrL1NvrbxUYbykLQ4Cv5XK0YCx5b4Hc
/X5t2z/ISQCKCy7qO5Egce4ormVl1O6miFdHtnBPveXfMn6K+GxUURst+1abYLJTRYkftY5HevyE
3ANv48sg+YHxraNvU5AWMtc1mYsdiUzjR/XjMijIB/s9bCichRR5D4UwRmDlj8qdqfGb90q5KeEq
vZfFBljclOu5DIlLOdW7kdekDWNA4kS/5zW5eny7R7i77q1j5HfCe0HueMBfHj2dROESMxF5x8r7
ZgYG2oEDuNfVWjlJx5+btRP15qWMV0oIkNMc+VJyDmckJEx6g6IOqb+lrA6iMSsbeQVLY9maPQWr
nzj1LlWlcq8MT8qD+17OGhXs48QhzbrKzNfbM7xbeu2oxCCFBfB5NSZGZsZ6G40HrKLaXW8IRsw4
e3iaQdWwXOlmtyPlCxAeujbVGfp9SLGRYDKhx+zCVYbPDJnuVAOzi6GbLcquQiAl54jqDPQzyIA+
BS1BTsUXvxhqobsU4vaGxErSN40TzeUzng0e8zurPQsGmQflB68QGT3/yoEe+twPO0e1WbyfDiF4
IpjQwFgNSXJO3Q7sI3QHS26EWyRSxKMN9s9YXEI1VAVnFYl2v6A5+YiDqxvDo9+ZFZijlpieERmk
1EbkuTZ5/UaZ6ZnZCRGQ9uWgqWdUQMt+ppLYvFG9L1mvJM8RpMROkXbOCjxNx2v1IBke/ktp+d5R
HjSdufgFnWWdVw8v9jPK8Szy0OJE/LTY0dB8D0jIoB5CmFTKwOY+hlKyB4OMTWWKivpTJUPxIMNi
cwvjaMAwCr225xM2z0XcjIWj6Xo7wIhvCCotBsiQANVt2O5L3vTMfskqJu9DyoO02vXOmnn1uQEH
vheLTiu+G+xY1Sr0I44lGcnqxbw50NioM1hLSPgqSn3owFtZDp8xYaFIZZjIR/BLSaX2jeAXaF74
GwWY8q59VtFsZ4pQrkvkDOyA/S81IBANDBTqfsNhEZdPDmh5rft4zPkjSoF2JTIqHpiz5fqX5T1h
SZfsyZqHdcgmcDXc7sGOE4nzwn4nbHTc3Sf336iAqziAjHYt0ctaETk8BcEVrXBbOdOG5wxhCBGZ
LY/jIHYd5PBGBJfm6263ArNdn8Zsq4q5RzzshPF4dQ3h1hEYRDvWwXOticafs0oWEGNIbPeN7jrw
xcMwveBJc/GC8bB8Ojj74PTquhnk0S0twyjlXj644mQzsto3Xx3la7cuUJfIkFY503Hsvs1kWKMh
WyKYSChOZT4gtPW8a54vwYAILqTOtn8/LLM8MCHz57gornV4flI9AN98TtHYZY+rygZJ7K4UVBJF
OXxjVTV+Vj2lb+p83iGQYcsHEGco81pE2NYaVq/I45ItJ1Ifvt5nYFu1slGjrM5fROepN+Q4JnKP
YoDdcAyEVv9IyLCmB4ug1jx5Uk969IzRPeRBWKHpz/yurK8qq648Iw9UxIbtaSYchY5XDgaxbs6a
Tim9HBW/IBT9jFH3vIBzay9+QBnls+cqFf6Lkju1MUp6jXDCycXpXP80slJBpXI80tWo1rcWMrys
/n1iu0PkO4XDiyLVu0erwLLH8Uf8V97aU392XYqG6FdFiD0kV4tNdK33D1ecvcthjh/g24r7YpQ5
4H6zcpGqbI1AsG2G8qhvKg4eFvNSDPRi54YSGc0+8n2t2QAbVe1TnMyKKSxKnuATUwC2Z+u1IDzT
xcX8bATpnC+FYmP21gJmUOHWxgUjz+4AAj0V8ZcvRNxOfwEzueeEXRpcU3xI8oVT8iN82IwVn42H
hywCLgz01ggxCyRZ6Mpw5oBOpwKi77kDubrH5wJqVWvtGSrslCkh6McTbnfV/y+Vs/9M914RlPlD
uVX7PVJw6Q68KrPidvCZgGa1gSUarsElSX74KuvBi9nkNLyFp9wCxMYUOT203nGrHaDDbRiYIFby
wcLLd/wQXUzRC2VS32dyOc6lmiP6kUzi6Hr8rJ0VNQEr8L9VUJWjHeExzg7wdcVWTcWhOJOcyjZM
nAzPr+r4WXZ8ukDhcp6/2iA1tGfGW0SHxTA8iRRglHmK2BW+FwpHVc7pTfAWc/xMoxXm7XCyMEKl
lo5u0R8wq1Amul8aOK0/C++LVQWaKDtYH7W5dAY3IeVtpJ4+DHY6Y8wnEy0lfAmdFhfoxbO3x8OH
Cn24T9mRmX3KeYzJnsxOL6sJVpGEJSO8VAC5CXva4NPDX9qfN/BD2Ma6hkF9D7MvwJ8YmFqdvYr7
8nwN31L2JiN0B6y/Yp4FsswejbDmisK02kQJ48y9vojPVyOfNws47QDbz4WeubKsTNjV3CET+iVv
/yzvtptMbMQXnKgeUktgX5DcNpqBWiSCU6irEIkIPCwpChFFrB67KXUvHgtTAZu3LTZbgeOUxDk8
uw/gbCg4/FwH2vKL0ANYBQyShwgMo0yyWX0VRXmtUD0mDRESS0UUqeyFn1ieY3JCWg6DXelgfLhG
G5Ngf1r/O0Rv2G40v2ihGfjlUYeop5ZBelVgi7pad8bufd+yVtdcXaK6fmkYGPYdlPWHeppCY2Uo
dTPqC948m5Lj8GOcRE8u9mZugHo5LyJX051PHAISzL+w4qrFUzcAguhpGoS2IIl2sJNovY5CyQOf
aSbzxvriDdt+1s2m/1FDikl/H5zvzr1kRrDHuvWL5KlAElTYzuzjOUMlXqWVqMZLrd3IOgZpqJSe
WbPvkoItC2xVjvUcThysUyM4TOM3bgTWM4VwS+U3eI/8tBGAvISbn88/q3nOwAay+YrdkivZzXWS
Nys64MshiFd6ICvRArZ7VbfkMxB1kBjiQmR4PAtVAKIG0sa4eOiur4VX3Mkd3Z5BgwA/N91fhIn2
iryY042ZRapM8N5+jqUA+/9N1QGVxGV1Ia1M5zbNuDgtFAHMZxWYbfBZQ5BOZSCqi/0zwoyTSSI7
N8POc4gDqkJzIlmpqq+jM/Cj+SH/kBxCNF47RuO1JG5XBFybLR/7c2EPl3TPByMzg2dxEety9/Fw
BUcPQ/XiggHIxv4/2fnS4TCyb2kc8LJ+cFY2dR+FGFxnVyaB8l97suQUDfCdLWrt8SYpann4q1hy
ccHTVlTLvRzPBvo/f2rBdxjUA3T999UGdbzrMw14FtEnbSzOq7VvOUOhBqC7fd/CYlldaWzkQ3Ud
7OnP3CR7v6Z/seA0TuywJeWWnSm/lt40WCRsSwoafoUalnsbsTbLKLl7CyJ5BjPnE4bbn+vgBd+G
9Nc8PZtIxd3fDbhS1rzlnX9BRfJozH52iaqCTx02WEkQgvfDRBtx0qHMxD3gsreUIV7t6nrdpsAd
xuMi/J955bvv0qOPAQTKFEV+LPBe82+xDLpQxc17Jrzz73rlw9bQwYK2NJRfgWilKOIOk93VqNRD
grVc9qfR1IHl6WJM8ovjwoF6YaaMpT9WmaJ7INEEWgsID1dNdVYlPv9V3H5jhFZg0BuU5X7y2rNE
aIK43c6MdBJITMW3As65Mh8FbkAt/E6IT+sJirHlKWS01BRpn9oTsAvAZ/0/oXTOUICQI2cT/DAb
7OBXhVgwIahsIzJXUknEiIvPKyvZlgsQnXCnPUnUzhatETKlxB3mum0qQ67U8M5xfL6ga5Rk7EUI
Ip1S939uOkxEvHfS9rbvcD13dxnbD2/ZGBnwfSk1U/DvGRqsSP4sOUhU1sFnGHYs3CCqSBo4oc6n
ueGkiNWDyt6iZou1bs+zoIpzK1MlPWlkiYBGntocYJlpUAI03NKjpZHMmOjYjL7CErwQ5oihp5AK
Zv/nrlDwI2vdPoLK6pNlLsquw0Vjoa/visuWrTTk+WCGeFBB8VU0kb1i51Brjiz8buVXq8iOq6ZA
81P2tkyveegwcg/98mGTrgQiIxe1Fs4R6POVwtp1NK4FjcKuAdQQaSg628csL71oA7AUr2P66WXc
AF9j/hc20Em9Pj6/MxgfhB4L5ADPvzBABCNtlQU87bsCOOcAbhxjGCWa586u+fKtZmuDR4MdkH0k
Q66s2+OCVOHUIOrXpe01nBV+vn1t8eBvupkVlwYe8E+KtWjRWn0hlWdKtC1yw3gJkKDCydJ/8Wh2
BPVguyAmxrjSVZPBd9PWOAkzlWDWGyl4OdrX0/a3qfls0FY78B1Elja7fIN8dw/fyVrl3EqNaEfP
PDwcQ1aZbhyCbhOkT2zqUCWPJ9R5BonFqumUde3D8CtYQo7Amf+ANVvRf6wMRrjtMM3AjdKDM/GI
vH3AKZjNjr21icKvIJ/IQNmZ1CbP9VhHbzkqTxoNfSBo0xob/udkIggIbUQT+Iei4TkTO2F0qBfn
Nw+sxZkiOrHzrZXdLHpXcHTm15CYRSDNg4jZrHVYle12pD6Xr7Bbisi4pARFt2u9ondN2XBCntxf
UduI3Yw0Is+HbpWZNRtrVEN5ECUAJSKFm9qS8IzXW/ax926mB/5m52rGL2x+Ijp8tLuaRlbtKOYs
PcQJ2K54KYiZyOHwU38C/Nk49wbBjw0ADSo06AM7zS++W7vwYMPqZPfoEnaqPEG1g9Mt15SxyytG
j64oXcoVDHWcWkcQYZYGQ7okmz4dfkuL8kqvtVdPqIIBHHRbAmxZS8mEuJdUkfnCpHF0G0dWKkHE
nvKSCReVodEYFNh6qiqBFpjoPoXu1Owc5Dkcd5sBkq4B4fghok/GoPmGNBSL/tK7y5D+V4JdZjsJ
XIohWMbVAz/YrcjdQRqT1xosdKWcs7CJJpr8LlBVBYkS+xL9tPuk0ceCIRo2xkg5oCEeGyudd0/T
K7HJ1JdzKiU5PkrdQJ4aihUGntHWqRs8VS7y7G2fnqCjp5WcAk7gEXGRovH9AafTDjMN+AUV+mWC
l1jnfjqey9FY5LCXmVrVAV4hLAIhoxlC93c49516ibNMxVagh/W4sHK3j8Veg+MUw5aafK58L8g9
nsVJS9MaIFYc7WT1/AGKnnZiG1BhBNvwUpWKuIJEx6D36NMvLWMhXLFBUVzhl9KMiet2m1cMGW5N
i/7VmmMatrBaoubR1lts8EqDgZfWzrz81IXuIvtjrGsEFmgSPg+aj6MzlbLy02fNfufoQnTpM20m
ZU/5hMTWPThEJ4GqGu0yAqxLjrtPgE9rYFajZ7BG1p1RYCSybs3BIyINuojYfsqlNcgnpyddeiCL
syot/Cd3+3vy5jJkmWwIlpAnZV1684lL5iag2I31OV+ojfCMr52x+x0obOlXvqh5W6kudtKrGgxE
1CQZG5ziDVOSIz4Jpa/NXdNWek5pfKy3nuyR/bY1sQGOE0jfCUekuj96n3W7laRXDTkh40M2hriG
sma4UkGLh4Fol+TB8tur050Wahw/kLBlLo8WIYTrgZw+tckf0MsHDc/a8ggeZDSd5NGLXJ50uQsz
u1s3u9yDSmliDahtRerJEatwf3F6+oRBH1gW+uAge4gg/VIrsusFAA0atLGP4JitGtCAD6PA1jCH
lZtAE0sN4ba909jF85KaPzDTara/juzLJGoD8Pphc40EN+KrdNOUXqePyMbFFmCWNMeJ8UTQ6kQV
c805ql3083Izj9nhSTfqw7GLQzUXuWlRoSyimR8++oRfvF55O2OStTj4YYoRqxz+kn+PU7x/13H2
cwn/pKZ9wFNLjCe5ZDHwG885pooOeEyQ2Qn3hoobc0OIR3AKkAIz6ZpBj5f7loU9LNgJSxNNhZcL
ueKNPKHfc5F428C5iP4fsLeBatjq+W9xP5eyvq4C3uyStfP9znoQCG2oJ6oCBWwfpcA2+l/w1+VQ
xKAJ5+Yuoo57MRMpblBtpf/IW9gaMWRw3sLC7I3BGNjfLl44rk59X/yyVuA8v4AzoM6HAXVaIqAZ
W7ZHaL4QFLG+lQ1o5+OOKrGo++2teSPMlUy+EhSmYeRh3ipeaTZxmOPpTFCmlNHuRHD7FjhAKfXE
Y4qIwQaFw8gohpURIj1jOORWej10X1aTM4c4SVxlq6nLXX8F5WtfIxW871glwlVnl9+U9GNVnzux
cxt9Nz7+8HTEk+cOzSuLZy8mjrkznBetVH0dWGDsJOuKgQkQKXXrV1r4En7KmyuK4pom52WnOZKk
Ov0dYTnjeuMrD9skM4/cWcZZioU9bMYYwuVTD0nafmYJJMD1zTWcufwxfcP2A4t5Cubn13wUzAlX
GKBudgCVsnNib6yZuot7IUHwC5POKJBKY1okpgRmWwBY+NuRHgjOgiIDnD/SeGr7ziwfo/kSn4vd
adh3H74EZqZu5NWFNPMH4eIwr3NQCNGX8qRHbVZ2K4e94LxbzMbbhYu1LW+WLKTtm3qB0f6c0Ovw
A/DFsRdMpjcDDvCqahEccQrPQeUAx01oBhRD62eDkDZeAiNwBHy+ppjM/pMABmwxwv4y6QzlybDK
ik6fEZjhdYjYEKwcDXb4xnNe8ihUf2V8lTS1Eht/x0Kxm7pxM6my/Mg9mzBk15neWib8q2LEimaV
5sAXpMP6MtdizsncukSN1D5BjVpc32mn8GTyDSE6MTB8RGmnhjKo36nSbDatfnObfjAZbPAR5zAL
i/mc287efU86E1S5Z+ECRxWf7W5n1QCd+q4Dr2y+4KgYXXQcHZOWvjq1KDRCTudcRWRS2A5TROBw
NVvmyc5qkLPtegvkFjYDPy8Q/eclNq7bwitKGmvRzK3qSIrTDdPSCXIunW9rMMnc+ZYaM0tWC/1k
qpMweR6mVOqbHvdXDQESLV1j3HXK3aUmQgsoD2Hg+1qLu7oLu+jFFp8DMao+AhmXlFRPdA9OvTxP
aFfVPvA00/g/TSm4hH3KPaF1kwASFlalKcFke9sBD6Ohb90z5GGFkFWEsygZ5I1SeO3LleckgHRE
Nr8fiq2aJjobKOF0uZiKMLVqKZPVvSG+1oLCIOXWVTih9eNpeDrn4yNpM0WdxrBsiJM37+v1a95L
+htwNFe7Mo5dlOKCKUAxC8r80pjHIx5POoRbmRd7+/6vUIklu+RQ1Hv8XZVLmX6uUE/MMrC2d9F8
nJqepgVlosbkBGNinVwwXp0KGPH9mH3nhZvz7PndoVQgWFBFbpQtF8A3+KfThzAuLYElPvYvkcT8
8n4/sfuyXgDT7tkijLuj4HXIuWcQzxq0kre8gou0C0vuEN2JrDhxDSLC9GgPqcTDujmtVikEGKJc
h7Payu8761VDseZpzHUjw6ngsX+2nCISeHmu88Imuhe5vR2eKRmHNQub6slA1gvTvNBhzgPfLIgf
sUNJz1j0lNH4c/f575gQvpzUNRu01ix70bvAXHi+8fWtFS3M/eoECntrCpFPGZDF1jVFHIoRwwnh
4Qwb5jgN8hsnp6vShmtBfdMCD7Djakob/3A6rkrThUqGgkRj/DZDKwj/OygSD4XpOAbbDtob++Iw
vQC2FYYWbB6weD0oFJ5K6R30yYGIvUOO+zBzOgjT2Oi39+1BrXup7pD5h31DYWU4rzdALceWyKO4
KbWMqym6XOnEXoiir1k6EPqXwnobi5b8biHnV5Ehnv0bGKqO2FcVeSUywpvY+vkn2O/7h1nyd4Cg
UWv0IOYxJJ4pzqtqeVsL0Bgs+OgDYnGQlVkZeV6J+oUhkZAUPjoW56My7M3Il1Ls15BLmK9XKmsi
gjObG/B2/a9yLd6lnwUHUqa5OLaa7rGu9tWo7AFJmHXBqOfj2Sjfdcx+3euT/SnZ2NP5YxBrPmSK
8xPl1mX+Zkfxy/XBni//CxEHz7sacj+ahYMfp726ju+6tFSEtVQS+/VmH15EbDfIp4rOBs5bgkNA
UwY2jE7f8lee3jizL9kdszsFbomrfpWVCIAD1Tg25STPAoJf8I5xD3v7S1iZpoaNoRmc7NJlABu9
5Yx56o5g1uSPH0m7xxf4Of7ywtRChGuyzw7OIl+HB71ooVr8NvmkB+MIjarBO/Ff/taVlx0ZPO3z
CVzZQLE7OxxHzhdiD0pd54K/6MysYPzFxA3YgzMAulLv9yPTf/JVyCpI9m+TuCRCxhSZlz69p1Yl
2flsN4xpSBF8SL6xH5m6bv46lv1MjyMV8jHcR5ECjg51PAGXyEt0KoqYxhAUJcpcJjVZEXah5/bM
KaKr1AWTloBL5D1SUBbed4W+HMaf7NtnZaaCg4zhtPyI1DrCePKIWZEHLi5AZ3bpK7tH7jkYBGLb
tlGSChy4xqvlSkvyPAfveZdxP3zoLg2P1NC1pYfcQryLesCQOxJ50JA4vKIcBIYgLf1sciNvHi4x
QNjB4lGNDSTeW14eD+Tub5DZN9JN5bBpHLM+oGhQc1Wj/Aarzt+t45XWm5JjV7dF2wwKUNOLjkcp
Ji0BSXxFMhijBuNu2kFqQSyF6jQMBCf9mvg+rUQPBefpWF2FuxlL3lb4Vs2oTMi+x8PRPxzJeZ1G
2neLxlPxJAyPQX2EgVny4l9/3Dm6TGHzUTwbwCQ411Yjai/QmzcqxYFIwAcPSwJYFuh5h9KjB/83
BQUlYE04lTRuTCTv1hVIFWRhq+JzYnQSg8ZQpE91C1AoM0eMGhYfDKk/x69eCcFSe0iK1UPTgPWZ
dsbvbmd7mv80K4/wlkhefKmMWOUUR9jxCOl4mf8ueTvps5i0u83dkw9lZYzk48VmG9WmXIgbDRT+
NgG0LPa7EEVQoT8/X0ZPLqzvB84OC6F89xkqPvFWeNK7meniap4jq4ZUMha5nwbv8FPzv3I26hei
MXkqP2O0npIl5A1dIH5uAA6oF+zMX7+YPjwNn6gMsgUse+uw5qmBBLGaewqjkKaFlESJqKqGkVkY
J0G2x8pxEn2/mwwh8r+W31bp+Dg8ulanpJ4Ivu2ljk6ZWnDI825AI8vpYyKa0WcmDPLQW9i0/FvK
cSQFbSAG/Z/1FygaIhh/dhUv4tcXNpembDElNayvyLWBIyj31swlbxKC5eVWncGDPaZOJUUD/Wgv
WMSj8h3M8D4/+oE0xCa4qumxVjAWuuYYycNSM5WOSgbmPfhlJZtlkztHlsSeLgDOFnJUYFv5tcQy
y4liZyrRy+vNBkD6Q21ATTMViFGBkKbjPgJdZUbfFw0lq5T6mk8YuvoTDPhxjbr3GYnf49yXDbVy
l3+rhlurx3nyQb0Y1bIEcBTUNulGPDOQtq2a5EARK1Yx3qALA1z/29E8LEPNJGe15ufNMB4ZjBas
gcppE9JbntN1Ab6rFZSb7RsY1hvvXFcKSwnKZTNcuEdDVCJ/V7+MCIIcf85xQ6iposthKsmAmoyN
m+c6lo35ysUFtMuD7SSLErpnE802yYDVvwpzhdjJC45ADYhRNkxjTQBmCWCQVhl3d7/HIcti2YsS
2b8ao98LY4af0N4wSwLkOJ9re3YmHS530x8RQ2ll43ZP1iE1L/O484fTleuZ3DR/6nmQX31j6+LK
xMD8Kptqzo7gGWhqKp/z3JscTet0tTxGhR4OGXGAQcOAvAwCrnrK4Ht32NV3A7bkK7X+5+nlfrel
LeNjMV8uqMtTFPQ27eSN+DRPg1MUCiM5wLDTxBk9HxlXMO0xo4YfLLEjVk6uKlgjr6ys1f2aeMrx
DVmS6GtAw7/p3oAfc+1d96a094oTBbJxzlt/ld9kr3iha2CRV83wlQwwWif54u4V1IsTGw6tc/nS
mgz2s16lbRIZgRBQcgGvFJe7uly0DLN21W3FVa2G9LkS/b0W3aR/cRCunaL2Q3wbfSabADA1hWvn
6UH0cpwT263C+yX/a0wPxc+Ues4oXtdvtl85yq0gf/EdHx89H7UMXLoAdGMgr3hGBnlCvxEDWJ9a
LF5p8RVq9YgPPA2e4s+TZLz0T6SStZMnqeMJRfn7LVIRPAFA4ZxDxB1iijFIqinpWbM3lyppYUqI
iZ4JBtDL2kDjppjcXChJghdB0cwvbtLhVcb/hRxuPoJ1EtPF53yxoKXqygKQ8k1DTFPi8BQ5l5M9
9SAzK3JFd+vNgxfJA2vYdRAjak5ce/I6WPiIHIwP+G3axaB06H4UAHpS00mxbxcbCyomlPMKG3Cf
3+zkbQ8fFlzr0diVcKm0Xe0dtxSaNMWozyPCbQu7b/0Zx9vOkqo+xWjGPXRWLIsxef9JYy2ednDF
EGWu6fztV5dRxXUvr0euZst/RjnSPHa33zH85RpZ/CrenjNKWmwxmuxh37PSpw5OMvF0MIabxSJI
GNnK019IClOOZsKeHfAcuRcx4tlVJtl2ugoMaF2tVEBR2rTh+ffR/0GaG1+j7DRlVLUf+Zl4paYa
vpa6uAxT7F3sRFx0p27mOSm9Xq8va7xSyx6eW7AY8rkLfPVPNr1ifSrRqFBxNETa+SpQTNOSf8dS
vBtJLmOyE2Mzr7c1yKXshmfZTbjwyaKccRAvnHXGAZhS87phDFG4EtHJgNv2VFeppRoWR+0TqNkt
wQhN8+2Z8co5hJjKcaEFyItNEaIwrli4Q6ytYNUpDXRz13ilbbz2bg6VIt7HvuXyoyK/f6ak4kCf
+z6Oxf3v3FU+EEa6wgUgCkFqBHPdQ638GPDE7C1nTCnr/prvR0BHWwTu0VSGL8MrXE9BN++KeHOM
uxw69rjR0bTorSMBPHBVc61VL6UMOiyShaj3w6MCHgdq0iGS2qrGd5llmDa2t3es8kjt6SgdGM1v
8+R4jh3nlLDAYMlICENms0b2VtLQsPcPDuZHRqfFi45wNtoQVbMzy8HzI2qZutlPqNautgOO0fYt
EJjADSfYAa99580xxyKVN5tJJWHkPdarnzO0LAKXLZfXjFousB2UXNRcWnzb/0HikHJk2GokObAE
p3zLZe78+SaMK0WHF9R9FBiks+MmK1bMzSBuJruPs8M+80p/tvAjqtw2fRiK29LMCOhRtk0XcLG/
V+TlVT/LVH7OAC3e8GzqAs2qCzZqmTPGgtxn7RaJCDYZSRK8p+lLUq5ue1cT1DdwHtZE6QqHomc+
RO3y48J2iD/HtAzkOQa70p31cNc13zq9ZZkK68heJQMQ3WU1K/r9rPwgLFSvk5lR3y9W7bAEjwE2
+bEV5MJVZcHERVIU1Wi/vfPj2uFB/ZBZgQWs1ChR+30qQ5GvAfKI2lZU6EVKaQfKeJkPffvRLBea
Bl0jWl3LfED3/n6J4yKKUaXtI+eJ1Jnp4Ulv/XxkXCtl6JomLMnjKmTjKz8Qd241eMZ2wl1YxYuW
lSXeRc5ZwNd5A+hpWb0y1AmlpBinj01Igj2FIRiLzZt1peXZDcTlmsGYGl6EKh/yT5B62ZEYhMbX
ZLhqSw5CoYeHinwDrhV54DljMc/hvI3lSQppZIWCsj1sxgEAbP7Jg3RfXqG7FpcA84rikz4BLGVO
SxNRt50ixrmjKddzxBknb+3eWDOJtVnv8TXrDbdwOkmlUqLsMP3wsizU71t9LUUihp5oCon0HseU
KUiJprtR9KFnAJpiNG9205Hp/XyKeO5rNVr93DTf92yaShwUqsedUburF3cDzUievEBM3fPypLHM
i8s3p5FTp+BpvbQq4We9i+ppgoGYtYO6iBqS2NMjrfZiWPMLVeH0WNbmjTLha7D7hL0Khuqg36nD
NknORnemygEjtrn8zRbTaKoDn7LJAb6ir8GsS0CR/JPMWSNLC0l0XwdTUx8JnrDRXz6RGBAqSSPr
gQsguxsxwE8nx1U9DIXEHdn6qaPfLW0sjJc7SpNHfARKh86gO/M12a76u0QZ3gbmUkg48jeZiNc8
taBx/3dL1Ib18bGkGNk4++8q82rqPrN99/7DxfjdtRkb3j60HPT6325k3GHGRZGj3SHJqChXmadR
p1GlPyvxHruP3iIOaelWLbhpoxDUDlLeENJdM2zxCLcdV7Lf9GwQp8wR/n42nY16XVMa7KivUYaQ
S+G7kou7PFvbdhIqlZPgt0/weygfnSg2y51up40bDfiRmYgNKYuVr8xSKYycEoowPgXdadelWsZZ
AKC5djFjE8Fe72ER0aDdCsmA8hhj2L88mFsMLqXDDuFk+cH+5RecLhWyTC3TpOzHinOE9SOmbjRV
68ARniUYYTSMpKOf07/63g4UsJRrNX3wuvMksAYtkrUsngSUNbLdqQSrd0I8aFvTlNT741Cq4r72
Aa7fR7KCDEzVXRcE7MxVKcLsCwanhANDhXx5rIiDG6RBFr+e0Owrt3+ZWx/qCGw0ZK2sWYvdarBH
06t+GVEegnc6Ua1WKkRrV7cAVWOYa/HGgEDTIAPZUqVnwmZ3HvGoKjv+i0H+pBcpEezO1e/OoQiC
koi9iSkfhl4XA6UwXQZs6jnV8ki36xno/sqSYQqP7DRTeePtF5If9CqyT6/VpxysSorIU76FcK6N
y8DjH8iDBDMdf+MqouXNTJ/ZBGxZrP6l3xS/m129uOunbQXyekYMiyj1PWpcE3u3jUd4ZVrGqhXX
RIx7V66CokvbLqHBfkiXOTYYUh1NDPBnRMDK65KorXSXzWUF58pzUYDjmT0FkOrA9AeY4YYdLam4
hHwep/ydSxkbrCz35sbIM4ZKF6/oM8bwuRNcQooNotRgp/+xmNAvrUNzlFJB1uHyTxSnRnkezPAJ
E4PRk2S97rXYKanSEb8MNmf7W0mFSId8r1sysTke3wXh7shKO6RjGCSsbdmNvgJ5BgUeGJnXugj6
RSXbVNdu15QuMpjPqMW7u5tGuK46KMf8I2H/OyoOW9x17HQPoyuEYVZ+froBWDlb+BT/uqZ/VuHE
jjyTFOWSHCqmTJ3WPcVPVx0hmM4KLUucXg1n4xhhAlDeppU1RExKZxfmH1SkuAbGCuAdhOW7En2O
jmJ2KDydwExaSbBDOy54eorV3u04atg1D9FtqMaMbfDlCgwPpBY1Mf8PvZjVXaFpnn2WLBHll8rF
QPvr7U1x3j4/JixjQwgkKf5NgboxqXJIHXKejhNoUeWQG3PdhvnB1I7lHUQUX+LtN0s6UaUbFJIs
dDPM5hAvB/xobhg6lc66qfCXJCq1616EzvTBWiKlxqzqpPP8dpVynTuZ4ndcwhPgZUlSDDBR/8F5
n3GxpVZj1DODMybuux4HLVKIyZzYZGWwalapAgGm6s2YDT7U4Wt1k+XrqwxU+lRQKVgv2MadAyAG
+OkAB4oegnldWe5ScA83IV4G9V7A16sJMPTuHcVHV4SZZ2VTL/kp6JDlBn2UPzMqJDievDzvH78y
TdbxatoZ8GC+/hjg2gelGyzMbqdF7Vmz94VvwuUHQeUN9zoqK6fQaf3gB/594JuZgzvQekWoh83v
i21m/PClRTU9Znhgf9exrEY/FlQLqR0CxtRdINe2d9WSr/aVkaC/e/yR8InNqa6gktBPTYf0l6be
ADlN2iIps6d8h+pN9qiSZttsuHPdsbZ0ivObm2ydRAo1S2Slnb1PFtGnoDFF4MkqTxeoU0GVaM4q
PmNGEb/+AOo1wZCgr9xR99nf+vdtTS9Bh+nuIDUmoncSyfNNlztl70RZBDehIlmSbRRaZHt8vo8w
dE6PRCqFgYqOiwwurQACs981xnJT6WF1zUMF1wunu9ln+3FMI0JsJCKs5UxjnBlLICJLoMzYxI3n
aAWwnMkhNMAg8LMJf5cxfm5iuCjV3pI4NA/hxz45U+vTyJpWUDmIG/qCUWfQk4ouvmEhslXO/OYs
D6iWPTRaBJ6pbNx0Vn1dWl0a3ZfrBLcZ10f/nnYnLS47a5lk6h9HdhAnRvwZHs4VUTEUIwJek5tt
qWJXqYq8pA9pi2LsaZPYg0hGI8Chvy5gy97a1yVoTWeTe2o6ncpKjdkJ+/XBJGZrPI7NeVhtdr7z
U2HEqsI9eTPWjQAJQgMPILYgvO0d6xFru6ly7ee0JTUOX3Lh9PgMLM2xLhrXLM7xeVfT5WC7546+
GNFYarJ9kwygIAZSW5d3/ggxC1UN2Tqb5OIP83GnORe13068Pm15So97KqeUHJVY+4D8JwqqOWRW
bWksUjzefHMgIq2KSzB+bQO7f3wRt5WAa9t392QZMXjnkQK9jvazq5M2WxFJ9wTlk0m4umll5ZXz
zP98HfruzRUqrDpmKMz4olpXI93tr70g5t4LGXJtw9lyFkSkWfubW9Q3WY15JjSuhKV8ND8yXPnS
EBREcJOZAs2uZQ5GC+gdRYjgbkTFv0UQyTRhOmVtX3Shs8UfnbUVcCwrx3v2+QN6SnF2v3nx/2qi
u2vc/bmCku7SWZ8qgjQ8lBUlDwUzfdOvxTZ9+5Clr1LezEoGiS0crGFLZdrCStw4DplOMxLmW8n7
3yqsFv1Eeb8DZoCcxb7TLLE0cInPGxJzX+NoubnhJp8AYLXeNooicfMO+zDtWY2N6aENoQnBdOG5
YEyFGyl2ML0qQoEt4Xe1B5ko/wrUgk1lPTMpZvTomn4tvUBwfeH1wKNiA6SazwDZDG7WpyfeMElj
HzofYHFdP40Kfel0hgqXoT6xYyTLW7Nkt1NbxljV6fRjfBG0mIMc4jnOihZ0Mem5nqs0fPgjSYBt
YPX8IVVJgFCGgLwdIEeSIEGRZKUIRiWFxbFs2wTZEykJBmCMvdud1IZB15DLLDbg3tDM+S47qnVd
AqY10joT08U/vp7rVuCjIvGiWrgXQ/Db6vjGddjwfW+vbbdrI4FsXqstPKhBVmWonF/23kO7ab4p
QMhz2cigRi/cxjR8KXgmmKFizM0Tw0GDTOzLiGcxqFYEpDxagSrF9ZDy07HHH4pgDi533fBxC3I3
uJteKxwUzV1ZWZV6yJzZh2ZNG1u2o55qKxlZpS5S6ipgi22Tcv955PJX8Wb5snaS1VtRoqOFtpTQ
NBS5Ev09wd5R4/AKKDJEKb0BQBDhdyX7oJM4HzA8qLWSOp41K3ISnh3+/AqVJybg4juZTm6UjfjQ
k/5NMT3Iu1Gj9jodA0u9IeaPRYkbOW2vTepTkoEaf9v/S8J4gXDKextJjtXsU3UKRFAbFH/sCebi
eEV3WHHm0kPMF5EvYoYlhJn4UyMTX1ZRMytcn5uGdfYKlVTdW3pI59YFIkFstMy/ZfBAU3giBn1l
mJSgEPp6mWTk7r6rZJ0m4efk2IxuoQQ/X+MlvzmKxg2UmLB1nkzMo1GWP74Hs9TdYHb1STyAaMKJ
M37v8t9WDxY53H9r+E7O5EuPzPQdtVdP/XRQ/scTwx5njJAU2WqbxQPlbnLyOVAb2fwhFUJvjDbj
J6FQ+CRdilQNZIACg16nGBKOu6iWz9u+4O3TC2aDSH4cz0AJw0djyMIfPIjSfZ0BmXftw1T7KZ4O
75WCXAOUlyvVwMQnhn9siJ9vvxLgbYmHISAQTFxHP/hry7zIHmQnOaPxa9+siPjD+ACNMdG1aN8C
8URcA+4rv23/AhEYnop8J1zkNN4uGUpEjYXYLgN9PAG/dsNMCX6ZVfrMzDNPtY6KjWd7Sz4iqN0+
gaE3iDT6wGTaQUoCv1LUDNPW4M+sf7edxg7BGZVGMx0MPgrctIKVCw3cRICq05MYPRhs9dYbl/Mg
QVhEDylZ/MpX4k8DpoEQKvhF67ssAQToXN34gqbjKW2/ZMUjtJofaJ/THbNxkOnY72S7jQh8h368
st0ChRFhK6WuFvwnnTzSndygbaDDH5hPQqInsAeurz+WpSI+Wik6IEvgk+Azqe4+T/p5hfvKd6ZI
cM+2Y/c6jciLlZh4AU7pCFkJK4B2zkXcJ/t0lqiLgglvkFnrAeYS8Hgg86/ASQi6bPUcx0UuLaSN
9+QqVNsKWxfylFtYlMp4sR7O060d9s3FXSci/RoEyYs0gRlNqCfMCsd6JfcPvhsvEdKbqnXRxDDL
Dd7YNk+a/xOy4Zs+86n8IlgxD89q0ovpbLIE+4l9lOA4SV6Z5V/h8BP3HWEJuc2/6VBTSWCaQwFI
mfLKhrFMuLBtjADaQ5yoHQ0JUhhH+/0q0lsxfCDxQ26v2rxmsC2zkqeH7JpxeL8U+6M14dUzNDg8
mYwlx8AqcFlnS/Dn/iqS+Hl0tWwCK1eZOkZQ+gb1XPw/+yUjfrIhp0IvsxfUb+Ka2zJhCW298ubf
5MP63hAD6YSPPSZdPtACUnKcONByLHd7bgWaqc92cwqe6esGexRsIdR2iOR/7qSFBrPDqYCaLZVP
EJUoWaKcsZunTIE7ng5wQeZwwaeZ/YUulbeLiZ6fHvhNoTduETyYM442FL7BoxgHZRxFhkAT/BMC
TUVK1VBEvb4uVGTRWyLwRSn9sx1J8CAnQ7OS4nK5zjOJeeGZkmp06FNzXZuvHGc3WlnV86mWh1j/
AICRw0WqB3zJtrhIPE0pOrwLkmPC5IrBVZX3YWMXhTuYA7hjvR2StLjw+Z1YWBr8lIvkFke1SIU/
ubmoN4uzRqyQLyevn5kTkEpAWwmXcRi0rjzDT8IaKXoVXFS2Nhr/9sriiDGpHACX/HGle5Gtfue1
j8LTAiDZfuPgC79QHsdxiwm3r11wD4yNM+JWyrQncyj1VD5s+KB1Bkxyd7ZhzSo9BBj5g1y3KBhQ
yvGLwPkW67yibLmwNq/KWnf9CWaJgZ6XAsZapF02o+Huq8s284PTfOPHhZhRbSnW6ruHzMZRzQK1
e6WCzHRbBJvuv7ppegp7IZv3kO/EEjSxpfBM+JnQd15rS5A1TFw5fENbCIdu//ZE8xQVD5svQeea
BrV5IcWvZUDdiCph9CAMaF0GZWAebVj67gboYP1ugJTFnQFQig3PT2GuOVpzYCqN7Sqt8cTtLpg4
cvYEboesYdumWZU/qiDquqCCsRAS9+ZDhmm/3n+oC46V/jHN9DjoJsUSDtscrTmSJMcS1U1fmnBS
xo8YeiUqHUdw+9fTbMj60TZzMXOsz1rkxU2KSc4EFK7rjtJJpOj2maE1f1pyazKTclsEsfrMQKYB
R75N+Z+ZXfzpAvTcy8fug7S4EPvFKQI38w6d/Stmgu+oR/6PyMOjNV1rpo2OguqLTdpSQjKBya5b
EZ9jJXeAnATrUwd5Ws+hJ6EQRtM82oe52JXAQ2idaUHjtwBnMoRYk9cI7zbxfyimPHKcWoyM1JLh
gOMOaTDZX/up/UclfWOjxHvYTH7XwfUhQFc6fUPEFJI4IdMVqOag0AdhS4+7SbEe6Lo+9fyUHPJT
sqeaPVha9Hxmf8yAdNqhBozRtiAaOQ+OxBO8MCqwDE/jkep50E/TOEgbsZA2f30dIpw/lfWk6n7y
thh58uis7HhvWyPe6qe76C8C8A19dfk+INe4dD1pwIkW/usMpJ0XTXe3rJ/lQOGscBZR1VUpyg+/
7PdEhUUnxFl9z2kM5x6hASKagAz87G85D0L/9l2LTCsiDcKCVdgQmm+tTLaE6WJEOjraSau0lUVM
cxKE/Z2Q8xjc74MbuPc6zp1ypr5DrmZ2xCBk1dQFlaIwckvoqaPvKrWFd9lituuGLgpharBOBKuA
vaKeJNin+Xy+575xXKbHD1TWvbEEzhODdEF9kU0XxjKJGnpUAc3oeeUZTrY6vtBlWoAOsWgE9q+7
XKsab7cV1yaL0u+8jQGMtPy/CsWCVLKjPAq8ybWriAJwh2S+hh2Jbeink3MazyU6HHd5W4wnvBb+
bD5kGZVcL4m6fDLaqnAO230TAgLU6rqaZD1VuCyHEcObKttSac+WQIqBujlG6k7WTjxQ237gdGEk
yAtqUJTAv6pcmAbkT+1YefGo7yEG6G8YIZ1IbmGfco3a8+VrcVnpEbrRcDDpHy1+bXmo14RrXobU
2A+Qfv1pBfTPpAOQ5h9pUkkaoTgoNUcbYua1ecSFZhGCniGI0wBRV88Xg+GCsWQ1NcvCqj/JiLQ7
loSYsO9OWZCh7Cf4e5rO8NoTbigFxFFpaRBZC9XCKuPaOaWuBX8O8osmeXR9NtWR3WLUPZG4BxNw
TwTurMTUlq7GYjvBqsbN9XXMNNdZWX/n1NeMQgM/EzwRoTMq8ZiTgxO572REhTVv8PBJwjd00Pqc
ePuNNy84Qg4zgcGRyinNB+vitgee5nAdYheu4913AyflhWzVwzIBPEb/BtRsCJWDrOaM8nCT1/vX
Vfrmgf2M73U5LUbCHjvUIIpD21E0dkDoqyIZW6C8fH3jJlp2kWECHCAuF+HG9DXsXqGPB2xjPlzi
/BLfy66UgLwksMGo2eFWhC3Mh1mRFCChgpqcbCded4wgHbskkFQ2BsI+M0zCIVnHHzAWFqmnjsMF
JQpvTweaI7+Dxse4P6jg30zEdXtD9XO/PVxsswanEPr2VYMD3rGUxFuGP/kAn27Vo/an8LMAxsV8
7pVHj5JdG+/4Iye2AoDilwE4naDI5WsfYK+CZVdLLyz23tcG0ax1Ja3ShFmfTWL2vHBkO4Y5Jf8T
XJEbKByxoAQU1TkhdsuidqvKc/1fF5F+CZ0Vob10PtJl6PO2qiM7j+NJTAoymXgYIzEhPf5s6uTX
WtKsfxekI04q6yEiiDpZAOkGesX3k6neHei1rq9SLzOS/9HnKgUeq+pxqh6Y79L5WbyclMu8yQp4
KIcSNQ2dMnV5cRg2byDbmKhdrbnl7htW7HUjbjyHdaW4kXRL0Ofcj5BgPktQRuXR/UBRAClNAYRf
n+2Eu5RXPIt3CcGpo7FOt1gd5MjE+X4v4OhdJK59KY0XCVFAAMdNqRftQyN98LePRrnUle+7RDB2
hVziGAh+YNjIKdGU+oDeKXeZqlbg+tNMm0BGu/oqdKNrv+yStu0WZnJjh1fbH1XOyGyQBkFCkN4m
cqSgbsN4vu9ZnX1w5Fkudy8WuIkHCU9+RFt7tzb4ZMvkif5YcUimPhPYqNlhamJt7CmM54aW9URp
o+sruNterLdHp3jsi2Rl9WNfq76pZ4WYFkPSYd2z/ah+Ya298Dz+Sz96+7GurWZL4haZon1nvEMD
l9hhU5ckHqqh/c82DiYO48mRyvn4mBGyfnQ7asF4vMVgp0ddnfd1B1t+Lkji2dX8Xg326u5ah34Y
3ubfvOKuZALjc/KPvwXOV3fnf7vkQvDlR0sxuOKfWHJI+F6sfQfv1Tk1ESL3aGouGbV5NnvhoM9V
wisGXOHXj2Pv+zdssBCaWTnWtAmTt/jzcE166xDFaWLFBk2JgMPeV2JT32KZITdL/fCpeApLrAJc
G/yP7lL9K9p06woLAZexf3XgWntQd8c7MAfmjPhXG9C7P1UepsvvGMoafu8bD3mlniNmUvUQ8gHz
+3I/pC4vThJri+w81h8TqCYLastoMKdb7B5/e0f4OQD1yDRs82YBOsOTRVqUhFvtkpSfA8WwmiZA
5agjokXDj4jWVbQ7xTQY9N6mtw43v6UFdrp1+AE+GdTAX6O3C8Bd3ShgjzBzQ/PgoRDDwY/fHpdG
mIZxUsghJqiT9kEzL52Tf3P4Mg34eEF43AXISsmoSH/I0VjO+tV9qbvfS+zUD0iiGlN0lgcfuR8i
CnMrX0bx1TgMtSbjYzEboSxe0Niq5Qbw6crhUf5TAu9VDphmUmTL2Tx8kZU5yaCBobKvlGthfHvP
/HesyK1upaFlspBrdHXpOMCXnZfdi2JahYmLdxafMY9Gis02GxdR6r3vpjwtzNWtV2Daot1+5kli
ClSmeLKFLggw1eyryOKAUA8cMQmSbCvMwonScrPWDLUVM2AmOMzV9qklAz5G3m1rcNFlKPjM0ZOt
SWSIaFwqOz3uAbtc92I17PVV4d9OPMr8Y3124JEZHQtxpc7deQ6FGoL+peyAwlSWmJPas0KVzIEt
y/hB9OkmGQdVkBJ2VXWJJm42Rsw7ddU2sBbC7Qu7o3rgv8swfL+mEe9kyhw2C13CbsH+3pP8m5TK
u/kAnYmkpwEzbbB1KTLbOJaB+7hFX3uKP6nJPbZB6p16O9NbQ3sPsdJmjioUdgMxPilM9V1dpplg
w8KhNKyJJZRDoxoccRACmklpHDOtdqtGIRzgdDeehGuGspXL8t8XiDVM10GxqOlkE3DmrWGgnaUQ
1fs0mQGqFcrfdPPwFdPoxCmkFx9b/nuz/5PbIgYJWTGZFSdRj6d0IV6HVyXoenscSpWREwRnd2Rl
nwONxLuRH/ACJCXIXuwA4a9ytmsGGJ5C0IuSf+nXR8Igr1BjwVjIZnF4teEutlN9KGpnthU42+vd
OdKfcJSuOMGyjVqvpjs0BEReskn5Vu9kwGXghgwif4V59Dqmz+oLP0/rvV7LntArD4OdV0dWNcYR
tcHtHq932JGZl8l5yE7qb+C9YjZp389vsSBcOqYjy2GMzt09KWpYBNTfFMBZaY15RXNGSRNw1ATe
GTtvWa2Vv+C6JVoyRNZ6f19UnXPR1SgfFWicajG45onxoy03l92iA8/WLlcpiOCfnSap+r42886C
Yup+VrfMkwWBJMOvpJfZcLcRS05fCNzN8etSUO9VensHZy6Lctz4iEpozMzO4GRFdeRUYQ7TNN/z
eyx1eegC2O0pkV5xOgoja9yz3Qmf9/Zgventim9oxw22mCT5ewilovIz8sXcepSxx3dWPc6YP2LG
u9r55QSrY1zwHuPhFaVns5up8r/z9GSasDwJUgFp6QizS2lRd4bqk7U5/CMoVjz4HhaaSVZETZS8
L65OC1F9snwmAwpQPmjD4GFfNLWF1h/n3l8DMgRWdZou0wEUcGw3RL/bi/U6kjuMVDepQecLHnfZ
XHft9pdztLfjHVOdc++rRi6hZ8xIUR9jwfMhF4MVySMuBVOmOEiLdKWYUNNTmHcaxcxTY6b1aaZI
Dhfv0Jn48F/YrqHxlE9vF0wgYwMOuJJaYaDpd/W06Xaf8YfKzSiyPtpsVspZAoW8ZvsR/UXSf2hs
v/Pfz1jWX895nSqaNICZUbGMQCQ7T07jgV32OgU1HgoTZGfBcwRuhZwOLvLs6T0adJlPtUTCkQ3B
NgvcKUGvMLGvppXDQbqAH0y6EjXz5kxSoFJMeqUaz6PG4vUZWRdZJ7Uvr1/0IzRi/8nvphejzRca
1ItRBHlfFJNWZZD+CeF7nkYLfkXQd238xXCfLOR8T/pin20q8wVB3cEhg5yTfQnqo29YmtEhqfiT
q4r1cleDkjA71z1YXwyXq6MHtdZDGe+olFZ+J5Ct1I+5SVkXGdx7/b/ecnpyVViPoUXQT6cu7/ek
rVc1A8a+gkAxSns2Phrz2ipRNkHdkbYQSRRDV5WEiJP7KTTW5a46MugthdfA716NJj2RGA0PTsDL
pRoH13kovP88COVx07Aal6fcrXOt4JyaX1I6AVU9ROivGN+Xgskp63nBsS25q2IWBYRFzEcZXTv9
AfTK+/Y98Uh57T22xiTwGfFK7RA8RZNBlp65QEh0J8T4v2tPb3Iw6WNl82bk5zr4Lq8v08OWhMn6
C2udmR0VNXh37LysOx5WsWaafSHpIOPMUhRSYPO5A0QHCF2N4HxzSx9UHTF6h4Bv3pDls69Rh070
I7J63LIuQ8CXvBuqAOKfKosKQXhYQjKoZrs8ow2JjGmT13+3ZC7aNhVjuyNRVnl8R9726gGsnpYf
CA49MPVOGVwTicE8ZXQqXDtDVV6KU5jnEm0rM0ZRnXVENgSjxf4KG8MyC89X0J6JsdDxU/h0QFRC
zrj76p34B2AiD+lDwGlBw8ZPCwFsOuEQUhkTxfQdiV9hWDl+x2TW8L1px5A9F5Hycf0LEYACEYP5
ZivMoR+TQT8KTvaK0n+rSQt87U/D4jBA5ahoOG+Iw9xz4OmenA2XunkZyevr2v1MUMkPMwpS7u5Z
jREWDf5Bmo26ClMVCOPLzvAC/36aX2tWEoLPMTJMx/8VXknv4++JO78ySC0PmDa6wbe49RicU2He
crd4Pdg+lc0nPP9/e6lDLqWh+bamqfSkVbvEDVTQcm3x0gTKW3AcGEqD09XWcwuEpW2G4EcLpE18
epjoJIo4DXIuuR8pyAdTls2AB4gVDAp7vgKXoP36m0agtTVxluoBwtTxG64tzTKD1z2SiXNjgfX1
3prjvcCVQNBGRKoxkomTfmfQsin9ovgYkzrZkgXLWKMOo3XJve5HXsTbyfI+8K192mTutrvuH6aU
pgzvGewOMGyVZFK9gpH2qXt64Fi/drjoKxgxJXcPYrZj/9otxN07kbKIfR3vWo5PdbeHhzuzJ5k/
aWoYWlohRM4rLDFb6u5PNvmnQDKY7JDw97CYSVTg5hsYyGyWGvTClENLxaIEP6uUhco5fuB6knP0
bjzio/Y3GPEdbiDvHYOvNJdpfYRrjft9NJm88Bj0zFfWbFvwivxrIyKNncAOZbebpt8tXCxBNSS/
cwVJKp+k4APxvYD+IqHuv1vh9WkDgaGPkDZwj25PyvVkjHSBG/6/HlEs7nnaBvAVbvGwg/oP3py/
Ga7cWXYvFbQ+Eo+cHTiSLYgnhLkkYZ1gIiRKyKNveUS4nGz31gBACdejujA70cigZsCa234Q8Tih
JyBhKtCk4NdsSnn32ybdLeN9G8h7iTGx4sR2ZWh7qjJGJX3iKy7/yxkxKNmlwrO1KsI9HbzFCUgl
k8nHU5Z4FuwrJiyGU0ZIE3kZ6UsRuGth8tnmdv9O5Vx4/qysZuU3NP1rpihWGgSA+Sx3niKUgNci
878+qnWgRmEArd1YNQq7DeakfNCTy64zxuJT55H+oSkUuIGgqkdQ+6ZMs2+8sFAKbdvOwMwPYaut
VBfoJKZtLKxXQB+g6651FNC40OlmWVY2vnh/BKvnehDzLNdTQZTgRtGt9TrXNglNapczRPWgWzdA
R2ybh0OaOjbar2pydiK5/h6i6S0uEwHnSCsqSBiVxyWMC1GNUGrrDZlZyqbdkyIRKFbMJs5CNmQC
k+q5Ee7/3wAd2bArkfuPi4H9TOp2j6zSLonVpS2faxi1IDzj4P/MQICCSqooOXYdDZqHH9wdZSOF
D/XQDpg3+wmMPHb42gm919x0phbS/VF0ph3HPTtHIjPLTbXThXQ95bB9QUDWuRuNcV98Ab9JOBzw
hRgWvMtpVdytvFa+9AIu97kBCj6G0rtLOWRXeZNH+pLpZHo4+Kmt2+fCKjtzgXpWMNWZD7nah9Ez
TWhZcT5IGP5cmHUSNutcRggj1mhaZZk2UQjIoz1hcXTrYWrqGxczYqUiTGeTWMpaz7MJ8xZ8dUC8
p9T4ixVMV9WpZA33seyzyyIDznkpuDL57Y/qX2O4yzlbxaRiZKnZmcoC7ry87GwL/ctehw8fc3pZ
xT/PsxYT6WWV7/1Q3OP+KVFr8OyHr4yWvTQsHD7QpwZDODHMPDkZcXobiB5IHjQ6rpNKWeFUFWWs
NenG0HDFDlllIQi6KOaLvDSoF8q5LB6jw3qAAs9Mkwfi/bzJJLc1ymvwY2GWbHSNb/8JTayhZ0Dt
1hUzIg0XjBf0IIlEMaIrHadyB81fkF8kaFO7ksXwIiTpHbH96m9gkRRxYT01V6SK4+jHLDw2KEjZ
L5DUvzOubyWHRR7FdfALgP/4iQdbrCi2UN/s/qamMQh5NnyxD7McYvd9UTBybQDXEhgc4nDILiZ6
ptuolEZsgZBVW3BxsuB+ODbf7fD4I1J0KDW1372PQqRutHUJv6tJHJQMvHxu//zmGHg1hv0eZupr
HRJJRKPTlRhkUJAb46xUayxtqeGlY0pNFyC42tp+grZcjqnK4UD3Rs7a2B2cnmjbpnuijfJzZ1wO
BNhN+X97OZ4KhWIM42Q67cJQzMgfliS5BG4Uc9aTYXjk7Zhx5+5IpLY0huCkEsB4BYKyeuxTygae
mN1fKfblQhKFMPgbhCfaqmZFwQJkXdgEZ4dAQyVv/AttlzobhVP/5qQBLvqGtHJoTHtMR1yCL0az
QWXWhLHklfUqrNbphqwIHiZi8zTfGK2Td12zAvd3KbWQcWBlgqV1QBWsRHzlgeKznSWucMntEvyU
7l15wFDVcoYQQqCJJ2GQ7bDIiumpmmDUk+tNhOCNchEhOHgEKxNjcDoy174QKGCwx7S+9UrXte5k
ndZGII3wQ9reneUnqKeVjElpWK1H/6U2oEeCtwbw4+b2/eTqiCaCIo20C7Xp88FPPWfFwvHth+Ry
Jw6NUuq+YoT0Q7MTf0EahSeEEMTHlLExGTucHp/seHhtHLDoy95EBtrBcleJWTKCfXpkPQzWzOj7
BlarDWcVforL9rRgfy77NpRdlLt6WEy21EBveCGGk+aQoy2SKs+Mm4zj1sruUcj6YwOgAP1d13SV
AYESZZNTsByOwMb9ruNuRHFgkpm4ui5PMtSF5FTXTy+iy1ERK06Bnw2nkmm1cMtDbCQbVEAyPTd0
p4N6GKv0jFlNcploqcewQCckA1wp36EZ23Bf7CMbQ1EbJZ4yes5wwERpI1+0mJIXhmjeN8s5UISv
hcTxZWhOpuOKEnEvUeTd8mDePMRvxvVJKTqGpLR4htWSkrsjroeiyHuXkz4UjAL+g9gDaQBtNzlf
SMMSad/TAceLkQx+W1F68jZsO1JKMWjvFpUsuU02daU707W9wDJIV4B9PCtquT0Gb6LhSjc14KMN
eL78poXw4wfizLAUE2+22BxSyUOC+zD2r+j2uro7zKASCMGPAtF1bt3bTv6jUGCvNTQhAMyWzSCM
DMyIJdANZubY00I+/dtxsf0vvHibxAN/vNK+Hdlsm/wYoM8z6SfDm7wSzC6Bz01rdQd+sZL1FYPl
a1euyWWI/QXT4hOUuRbX6gYBeCosHTSic+OnlouMOq6lIB6DXjeFAjMgmieaW/9zULrpBV3EyFyW
wxOaI7yb0QykKmQm0m5CIiwaTYuwMBRpHkmXyvhI+CDYgiBqKuYfuz73FDe7fMNh8zGg+ba5k312
vcIwR9zWX4qaR1UDi85OjnoK43CeGKJVQKWmyVenqGuXjf/mHux7zw1/+Kr1oO/ARXIlI5QUme8q
Qsgj/c3vaYfiPdyfexLyvfwuiyKKsMVpi/P5/WKsSNyK6EMjHA8KRyY7t9nOCnLTzWKjzb745f6Q
mwDEMnk4GJCqk84naabsT1bGdbicGxzte0O+osoRFSjBbyRRNYKaX96TjyZroZc4hOZdzltGS8kL
cexrJuzCa+wDO2nFabOhDl2pt0VUpPa8yf6Igih06nJ1kawBuAMKVfgbRzHRyeTovZPiws+zA9Ru
WS/ik+apIYUM5PrwLWBnYqej2//CtdPD5bRzYOL1l60GIXoxjCAzuUKfkihrcHLtac5g7NPNPLs9
E0AjCxwUqnsz6xSNNc5z/43jBQCdANN+sCCkw9G/fTpHuFyM8o+LGeeFqET298wT/3r66HOtCMS6
eluOCIfIgI/zN/9iEbCdcjrZbaVHRwce+/jLRtyLS+WudC1yF3CA+fe//bnXRHT+ISYM8i9e9eU2
bzgTHaCOCMGdsRf5E9ySmnp3u0GuOx8mAS4DDU6Lo3T/jRFl3RmY+MTON/MatJI4ySDqLv+MLkDv
T6aF+lNUGd6AeqttDV/JYqrV/ocSGSg7MrHX/BCS25QzAisrHs6wso9Y+VX+K9oRshF/pNGi27q0
1pNa4NnnEFumWdtF9AWxlOsji7LRWqjmGMq+M1yl6N5LhYh4du1oseavZKdtxbIwK5MffLtewK4G
I9NURz0Y/wC+TTcqnrdhdMpJZX0xrrPvURxO9/Q5Bx/uHP8DSNgKmybC5y6X88zN4aeB8CYb3nAD
zHGeTMCQPgp1V/NwOQsflvnDzM0WVKDjIkIvBHE04+61e8NkEgTjNETcKvkmyvPU64+uqWpuiuuN
FeF8XTBYLTlNH/iXaKDIu0sia6nPgcSxSMkM6+CtuaAymrOjkNPO5UHGPrX9vsUOpRssKqDIfq1t
6fd18gF8QotgNS6aUxKkCoGfEIFL5TLhGsAGKFpxzzd/b291pXArVelrfY7ToZ01eOQWC2vChfdQ
bob4DcdGfnmtaCmrrdPunAuBjve/Wn1aJM8lFIVuqH9WnikZwZhomPWEBeoSRo5QznexBnQ0OjDA
pgrTz1RCrfWUeNPTyKB2350Twqg8Wm0vf+HHeHCH7muCIvitbQ6YDSm49bDgqHzZnY88SJksFmZz
+TuV23PkCWtByiRIJITXA55qzKaFe55r9tZg+2iAAz2W/OQfytB8HFjlY35hq3khRF+tlJbHcgW9
pWM/Wv14TGcSWPHMn6w7HGab+ETAQCKT/6LqPU2q9VgVhehNOd39pHjWThM5EwDEmOhktMAxFssu
pJt0nNLQnlKl/GU0uJWQmvWNZwgHAyXeLaOJW1guW+SEqVUuh2C2j3FmjoQa3I5TCoZIRi9s9one
HjmRDYoTy3LiZsAUtsP+UhTK08buN+P8gE1t+dnr2JZ4DnFCHtSBTpGFMJ3vGVGPJ4HtIX6bwirW
wnIP3jEokP/wqhhwkTUIMfJWK7I089y8ZLOo0+ofHizOb7kJzB4a2wTcRdIDjwFy1X2yWznCJ3Mk
QqRdn2/QJ71R/unAWuKNWdLI70tZjSv/edkFJHnMgpAkNOlaKEm14rI3fmluZD4oCcSK85fwPi4y
kCg96qRp7Oyo92zQYuwMwwRt6jnYcOJSUerZVGQ295/vT9zJS5bCnIJGUJI8pWp/4+XiotJ9CIxu
1vira/JH+uE2DV8kGY7h9qw7usoCoXV4GC8T0FIwdbNB0iuOl7fWDXXC7YBKCvAhUO/VTWFq2xqH
YhXItWcZRvdqEeWrdzDcRmtybNvY6WFxmrg8EPCfgvdrpy5OPzY1u+or6b+e9+f8IWkDwriO9ndg
SvU00TjWcKr04y3W/kC62O+ftH5K3P2gtpQgBuIi0WDOCia25uM03dXr5jHxCIJRYe6m654xiUQk
fIQ53/wKW9cnV61ahDVAlGskuO4Ndve6rkB22E2BFiPh52q1AcFnqDgf4nLM8lKjV3CCj2CZJaBs
JgeaWnb+QzYo4pV/DiUeYc+I+YJBRXbU+kVj3w8TLO60TylM8MOtOThcXtgQeEqEHYQ3oT/NoIZe
RkrNIlk1/3x/gyzN2s9LHm1IEAdMrGEp1+27AZOf5GRlsZ4dXaegoDvtk64WXZSEX7GvO2hRvxu7
AoQVXIctjQ7UURpdQEJt3GrCwS2b1xqyOuBM/fQxrm6VroIU/69J/SNhQ4KTmgLQmv4eDecAmXqn
LacEmT0Jcc5kPMgLtYi/KcNfi84KtT3DuB7jbgJmjXGe4rGE16q4t+e693xZJkQ77akCckp10Wqd
3Fa8XkbjTU0OTjzxDgAmvZQrP2sU2x59bHzfWCyTgAiwdpl3v/c2QPIXbz+KExyGiIQytpxHzWu+
jSpl6MISdN9QL1A63hTQxIfHaUlbNnDg21b4bpJwZ+THDbfvo/ykgreK+sSnX1GIV2g3NgU83hib
w9iZG3X9eYXT6TMRUrcAkqOh1ktIOlt79E0dfvlAhkTdLyJTJ07x/TSwcaqlS6+BmuxorAgr3ERd
n7PizNiLt5KeU1j9iKujVDUP0QELJYX78add8m7O8RFt4yMnAeKqApzQ/cHjHnwCHI+9vD9kpD+h
ooKbFYMttx79bQMsimQXqyEMYOwUXgr0f+lZ9N+OoSswavWopNuJzPHHIXbaEAswEPzGCcTyr2wG
v6SSDCdZlZ8nMlQ2hLwVOBQrcjzWuHWJrZm6S7OZLnlfhaCGMguquRPFUUzx+gTMLpm8KR1jSjzh
rM9M1n81PNX8CbHvJpf8f8g+QX3KTOgFbQAHHlZ4pKYf3/gXYNTYAJ9zDQlJUfo/QeAzIUs99XBf
r58u47VyT/qShWrSOnmRZ5V6eKYWKiXo81zKxNgtXGzpbidGTuKW+CrvIV6GJzKqUuI4Bl1xOgDa
B7VXmMo2UpjqSazBQvTJCJV9nmhVuSNCY6HOOGf1EEr2y3+OVqYWxTKj9Jq1mqWyI26qelPCXFy6
E+R5AxEl2JPg/TbBTuzxicRSSsRGWAeEBiR0u3hN29/T7OrCeAXZLeqfvXztQFUQI4LfORm3zVOE
ft6105sSYOnW3XZYg2WZ/x+JkospUzaF7g83O0s3BkHT7Ojv+2CpDM5fTuzFcnfC2TtCSHWjDW0V
uOBzK83qM/LeKf1S6xnL7pvKdcdJG78gDI63kOAxXxg0ksUjE1TZODcDNUotuxazrSv4IDqNcog9
RZBJstYbkRFfA8E4Qo1Bu53EHONGxrUZkzqMbvgWCSHsCZTwRRxGZo1gngjCZ3vjyLcjisVP0WeU
SEnUdP5BTorDCVwTchu+GY3vH63Ik2KcsQGrsIZC7e4kbUrICHgHtj3hfu4duF+vXPcmlMjtn9g8
rQdWzArjpTVOD+HOvBA82Y1tmgB1STSzcUNEkbztj12aiXuSIP9Bo0+F9r93q3D/zbd1kL/5H8k8
WWbhOM7w34niGG7TuvZT1i7xEwjUW7C8QptF3kMROEVzh1i/ic3g38JPb023SNt4iNfU1t3S1zOV
Jb6rEAcbbDfk1/eWUZZKayTl4cqRGBqnOkV9WAi2JN4gFfNSIjYYpWr5TtZZyd09NFEJbQ+itxLO
oqr6TRAJWzp0P5tJUgpt1GeQPJ0zqkQ6oi28Ppvui+ak7KNZt2LNbmHAomyXPd2yonwVAk4unjr4
SF8a7j+j4IqNHaiR/Olww1aIKPyLnEQ7Qjt0W1BGecRlC5M0aiBoU91C/yfABk49j/cm3AQMhBr5
KHy2JUwqs/qrC2oTTRHFNEY13sM+5zu0UioMlZmYPnC0+SfaWyi+YFwfXZfPsyJCEQFxZ48wYvEp
tb2xj9vSyXTh7GJlgoQwCosjDiazw0JQAjy9pUclYm8jOy217AVYiUApFK8YJRn4mvHCXheZfbim
aztats8aNL56E7DG1wGNjnTZw7ME8l1ue3b+S7app2SnJj9pWOo7Jw8MHCji0TA/ZUlMXfJAJ7em
I1OQloqPJ3NN85+2Ku94kLQxkqbQdafzfzx6/HY/KgiePrVtA/gRYJLCPS+Lu2/ezuwi3gp0TpzS
LoET+hVPBtkps2YUdR/M4E14dviDzGW5/pOkMBUbRbFDED5DIwweSvcIRg9Lz7kTWji0xN5icgjd
eDdPKVsUWozuBbBszQgwlH3u7tK4TuzLd3iq0ZZJGkUNYuQ0VwvOU5heakh/D0swRjlCFNcpjSq/
ka0Gde87OAhkUsUPWNVP54hi/1U/OXKeNaHscgl2KKxd/hkwl5Pgdi3sMzPTR9HT9shgikYsNRBe
BHLciyeqDXbEwl69nkTROdvDRmxwQZV+5VySCHCSD+VHp89/sH1tGNyXE8tUDarWJBZg35DzsPVS
eCVMWnFcmiDtdSpLY2TRFgCda4uJVD1XgigQZkY9szozdW0CGq77qPzTXhiCwhbPJDnVWQPFS5q9
UVkq+OMsJTPEH/rLx0RDzbuO+LJlwxZryAfEDIXEK5mSia96uk9rKD+4Aje6z+uNLUkoI0BXfbnA
3nakVNRdTH0j0b/+049oAYuyotNGnKnvH5tINScU+eaTTZd+iXj+ZmgXLcVpyXSaBIJgDYkX3vgW
Tsrjd66VNn8QFLizVqCwhguwV8tmWLjzIUgyhMcnks1cOw7nVkSI3+41437oHbDYFSwj+h5Zvquh
hpqxZzGbgDrtd30SuDwk6nTOS73LIfjx8NXHeY8YoZKxeQoBlIeKdzITep6eiPy9lcm57Lr7gaH2
ikw3arniYozfqG6Wec/NGubzxvbEIZAHGpM/shGMrTGH5pZWRVSPt+d6MWPWzddApEtAFUYKbbme
LWsSzMh2HUset+YxgUvq6Yb9/TjnUg2h8VeUcUKoaRbkavlCauVmYS8FbXM51KUHU22lwt7kGQz6
4YMfInQnMQQxLt00Yheoj2/TmwH8+9752ZZ7rvhlzK2pACQKIge+42JkL5VdW0gq03Uneam+3ZYr
uAOvaYT1j+5tY8dml+YyeFi4xma8ieeAKz58d/WS0gT673Gu4+05iG4P4JCmbYfbfbYwXnju4dTz
qIlW00ExQTx6rz2Rn7sNIvDYkPVU0xjkurYs/srSFc9A+bbz9TDv894jlO9gnz+hr3F/EZwXPVsc
KaP7V2SXuBmEvgPLDFaYhsaLi5rg4T3cxpvjaPbnmTxOKHaP5o1BK/6sfkgXrR6uImJKO4hOxvhE
cx4KuWbzdWqnlncYGYRQBDrP1ESJYsVh3ojn1wkHfX3pJwvZmRcJh4bk95hJSwXvIaGaKq14MFCG
TKTHE+6SdACiQPrajwOdPdGwpL93O9Dk1EMLZVcn2eDYxZTu1YO84ccGT5WnUdWI6UCmbMzcxkst
z5qljKKlawIF7loKtwmg4qKA5skDJGR2fdfn5RJ3pdShWWrkYmgzOThplD6nrAmjSMvPya9fi3+E
f/lKst3f4LU3EzO8U8rp7yP2wR37lv015su6Lwf71PfQJWy+1MSCOGNNByL5P/PGjtRO6daGV8XM
UOWUAEm3GxJqifPryY+9cvLmsTqlFVkEwVu3K7jBSHJ280mKuMZwojZ0sgc0bYy+R881cZ18E4Kj
Sn4V4z3FVTZnaplTelJbaE9jobUpG1E7dNeY4gltuE0e4iEHt15cXoZbgOhBSGqroItYAXOmMdh1
K3B6BAI0uMVT1dQxq6d15b//C2cA3/fayPcM53DbD2tvrjZU9llproReW0xMhjZkhS5K0Avz+YAs
heUwaTwgh18ltEMpoXTu+aRkrdYgkifFJG79ZwnooAFByJZW4EMXHrA3uXFE8Etjgcd4af+PvrEo
cQV09pAgb6TAQW3XhKfY+Ehqrv3nS65ZDrOuhvAy9LB8KdOW57HUpf3CRauS38d3c2JmtyuyX2F6
8/PeHdfokkR1cka6ubBkdYYRfvDrFvUyYJYLQtOhARaoc/F7vK4Q1BYpQUmsTumcfuu3hgZ+lKuC
usOdUTE1+1C+NHCSamPI8lBD2vmCBnIaQzKcZuqsXkes8+bfiXMoWJkWcIRRfi28ztp6yDRom4Da
1zo5kj8In3XiZGHQtmDaTi+U0zQUwaETPC7wnzItD2natPfUwQq7wjLFk1NbEI4STFmdG53aIe0B
PqDfL4bA9F5r7lGFE/aJAAAeHdg0QlRFo6vKoGVJTqBwpxHdnBI0TrGZEiOFDZMIbsQlESMNlJbf
zUlc7xOCxh2+ijySA8rk187nu9u+7fUc9lHa9j+5AG6ojdv3CC/PZDufqsOqK1eHJcz1zYyP0KTO
JMJ8UdYuIHy6w2++z3vsrTTXv9fJbHoKGay5n1GyMrH85Kh2OMORCOghevqgkXSZ33obCFXljyuL
2lyYPNsGt3fDDo6jQQ6T9LPIgr5yv7EDebBP8thZpJl3jq5OjAcCRM6xoDLhgy7M42ZzZalead05
e7V0Xx2Ks/jydC/bzN5aD0WgT/W4jtDl/4yUyAE38hY0H4FcpNFzrxB7fTwseLnYrKLA+U4MSuTD
3vGDsirtSezEnzvA4hynvJbY2EQTMGl8HDm57Cml1LJ7B/N1HNnMJ+6lP35j69elGJj+JVzfwcC1
7W3Zyw2XPZ0mULN+bxKBEFZEqc2imW21CGuXUSQhCfmF/bkWOVEaCtCt5bz23s/H48pQgwL7f3sd
tVPEbfRbb5ZKVAvulJICLzkRXBLVR6QJ0sgCF+rRH/JBwQQ9OuFWazVus2tfsulZZ7BxKjdIET4Z
WXRItFwtoGg/tviqQ4GF07beMrn1w9ttw8gIsdqG4imQ/IvQrgl63sKjtkt9BxDKSv7yRUHv1WS3
ckk1AbLtYttPekhNEfSA2lfKOWn2e8QFlEtYBseVBpJ0pDZH+U97ljV7VyDoYgHIfFoq+naplIoi
/Mdir/g9TMUo665ikxV8bL/3+aNE2RKyDDz3NSSxXCNElREdBCEGPzlLidlChNEOnuwL1wpEg2vT
qIxijKK5BGWd4vVE6Zwj4cMsP711ZddLmbDrI8s+Yd7W9xiIzvghiSygbxJtVcr7q/NaeVXb9C5Y
BNuDjn5oRt0e6C9P7uEaWW2fI02u82Jlc+tWbo+Oufi0MreO5iXdfrnAPM2UUGpn8eQ+rNW7Hm9d
WRE9B95sJ8gdtOYu2/o3TV2NOLc25KCOOM4I4bVNlOdOsy9I+mfWcef+KdOR0Tk2itgjJnV1MG/I
NVdrMHgTWdXMnzFH7ccBMZ1nAMTh1o/IQRKdH6gCSb0FPQ8v3PXuT/1yjBR3WWxTsknRwBw5Zd8Q
uBeNiLg7F0kv2gP/DB06Q683nzUKELbBjeHou6h8MW7tOHwfl96W/CpW1BSTyGGDmDRBVlXv7Gjp
3kY3xWHtkAqGi9umP/NPyKQptpkPVKutILQ7x5Erl31bMs/0yyIWlaQl8zPEITAsTXDX/+QpVplj
2CWnmtJtAw0WMIn6xLjP84ixd+3QOLm1v38/XUDtL9SLXeq1e3lOwmRDKU+4W4EJKvqM6UwHj34g
XOgdS7EIJzF7joWLvi77yAWzys0eJNg1zRiXCJABEPCoYCMQlYwYLI4JnPlNA5IaNnJCsvrhVAcd
gKT0dQeSVFBxHRRcink1AIlHNVOWw/rKrF3qYn8u4uZQWzgQFOU+9X9OTRGtHvT5yceLcDGGCoSF
9o4M1K21FYFvIT3i+QVQKlZSl//i2XUpjldZeLbFfc4uMs+0UzLMfaoEMj7cX8l/xjGY8DMuGesB
wN5ZahUzJqb5LUfUqIisrkQ6FwzdiCryIIhBJeVL3gMDxaPr4pfPMLnOOU/mayeGBQK3SN3+SnbZ
tUO2/LARYr1ysVEGChJuogpGkeZ393H8wgSNv3U8ocHM5Bl37lF13VoWc9MlNHg+WetBQZYWCaBO
nJa0Ed3V5W5kAwmNvltqsaLC4cQu9ZJPx2MLgpy0w303DAiEK9gymn3XkLAD6aRJB7Uu3eJ8ZA8v
LoFmLfdrPDaoW+9d1EVm1kRvX+rJ0k+ntdwgs8HOuaKcFgpFDr3+acNeOC8ZQMgD7nTNV09yi44L
rKrWAF/Gjw/XyyPo25fPcss9lVFh+cIeqN0R94VjTl3KtVBgI+Hk2Ju8rfpJJSlseiIE5AYhr6HQ
jZ+URVWfRGcL2dH45e3BfGSAmbk2Gy2JQcV2G3OOhPz0q6dpjX8Ks1lTR7z9uxAWnx6UAx9B1i7Z
JmArwVAH/FAkjYg6D2ytT17G/LPnxgruxA1i7XgdTV2XQ+6Z3r16ChMmBCqBHH29FmY0z6F5ST4q
pXIQZq1zi4GFdiErnBXDMqGgNPZ2qVEJeNNDCMeDiAB8LW5ErgK/yyew0J2lvesd3fSS4tFdXXKm
HPGIrRzpi7NPTeUyNzR6t5z8q8lKmm+nVzHibyRpH2GEzTzJ8TP5y2JP93UhAuBDQf2vReakgDBk
q6feGrdRFY9INRuVP4V8c5iZYjZWdcaRLHuEjTtO3AXR2WYtlsVVwAS+cKUzBlaWzfkQUnjhkUL6
9IRg+0xbQINCsyc7Gc9t0d1n/nZIwyvxcR2y62e7kGbPJ3gSJpeiAnoetxjzHHDalkiVnGXhUaaa
sXTqsfFrYvjgs+mpthsyHbxrQH+n5k7JRt2EheO9iad/tq067fEXEe4Wo8yv36JYN8Jg3Dlnbqku
+1W4uQrk8inEN4N7LQh8yGL8j9NZ3tR2Q/Q0OVVmcIg5HRVg6LDQDSIxIlGSqtQXhsRJmN6fwtgh
KQmm1cGhk9mDa3P7QoMVOeKUnZLAjjnhU8CYPY5uB0nd8/5sSiy9mBeZKTmMntkFSFAlEnk/YfoO
DVIbGle6xIcwXpPNBW3RAmcLKwRTBp2Kz2UvMMKjA8oZO17ltqLMpN1pFtNG92dJF1O8+XhscMEE
TD9+QEh1e4HvdrBB+XglePCHd1M1JsvMM+H4eHOxyqjaXvkNCww0g0DQhvivUZC2nvwlM1t25i8c
sSbhA0uknjHD5bTbzP9470cgR76As3Cyfo2bTzhpKNIs1dDUqxZbvSgdBlamylst9wwHscEEvGQ6
zh7mVZWGzBzJ1rSThLH0ne4EOlsPfYp1u+ygo647Fevxvna3k9uLHrLvZXWGBBtAz/mYmuKLWINj
QJZnmPnD41Zxix/DhxkWs+p4lNBQF7ETFhL5c8QjzYE++x2Lou7rkyMuQg3OSsRT2QIBE8wloFXO
pakZnG2n6FWZWUFhq9vr4WigVPRByb4As0xeHC/5WVpCWh/jZVoFDT673InkMB/p8HJ5gqchfw4v
P457MJHMCkIhEITQU+haIQ4Y2l3bdWpMYpGpU06WYuDZmV/BdOhJTstgdUewhXir2NDPPeJ2BKe0
WXgBO6AitL8+t/ZvRasomyZwb8D0IxMr49uSFfQuH2NgC1K4kGT2F6N22vory9U32s/nv6KF6rNC
g8fGMZOmN48cVdoDl02d0EWxpmKXuw9dkUWo8RMX8/41zp0KGViWDDSlDdEJQHVwVribW4R8bhsB
1SyymlVe+UmCuPkXCAjqkM1mSSec5g80OWSamcAyRJ41bjqhaVhneEVU337pdSDO5FDmS95B5urT
xhTWHyYUndhQ5G0aYuW9Czx2C86EkcNeQKQkfR5oE16khH2tMIljNzUkHGCUNOAsnFuuFdywSukb
39Edz6wuQVChsWFMF33Vmpa4ZZ/QfmptvB/Nq6BEjULTurGbjY3u5VIK7LU9arXXw9f6O8/IUF3G
KwNQdGgjJvkPl//ozv+qJHH1QewSlUY5t066dXdEuJBunYpaPnjniZ549vOfQIvlo7bgwaBzclN6
PyohjSRCeqGlSNdJcTgKZy2pxZVH58WWoA6hldvCQOPT+P6xJqNf5hJTDIvt63x1Pto5D/Y7xlep
myA7GhauPBmpneChzqL3odWyq9wYBc9HxSza/zWXkNEB65xEsAY0skERV12AK+u9U7kYDmdC50y5
QxpkMKeqLmQGg40LzGI4YQS9c8d11XKsB+T7rUyFLp49VC3KfZ0Rah6szMPbSvxZTPuutI3kFSmq
tBHBpC29hkg4EWeUOmynRc6HwlhEeEC2CoIInPjrTrow/0m0j5UzyaMW38KV77dXkN0fXdc9Vrim
RuBx9DX3TV56mhLmwBDwmQcLW83l8J2mfwpsQlvNV5XBSL1pWVF3NcZxaF+5Yfghq78SGCIq+sRj
rBFBRtYoLQqvo/bXRMPS9uKH2XWZKPiedj/Ogu0RPCoJ+jNJ8m7oI6fC/fEgyMpPm1Hmjzw53pSl
Yukkr+JJcz4anRnGZJEHmZ1qO7sbYWY2PrBPbTK2K+RqKuZ+/GMbNUBQ93eP7yepOesmdVowyi7V
P+hBXTQk4rwsokcSKKewZKdL59KKPlrBjfGdGnzGqgVq1++Px8wIFwgDXWO+qoTqsl3CPvzSoowQ
TA08HpCpxGZG+/fAZ09+xJHtKz2OnOyg829pCYx8KJGYfpMbEYjSs/pX4Mo1hK/UgHMaqvdeJ6JD
cHtmjhz7ug8RTkh4MKWLlD07CphASoiJKvNyfmPeumX7o+0kXJ8WvKDTwseDkN42ZDctLikg+Ge9
lTrcUnLSx7o3UB3tiFAfoq0xTGA44WSgvt9c9s1WiXGWXJcvD9rD8+p7iiQx+d4P9CiVEzTXsWF4
rGvcssOCLVj85M/sGXXePE5IGFfOarawIIKi7gvSrbA+u6l8bCPQgB7Waniu4V6KZugU1QwByCsV
KvP9QSHcU5VABu6rVkF6E4JhS1TeycsVKhhvIbRDCTLPhwBSjlg0n2HjpeLmZVsx7/cOfUBasNwe
ZxfYljwZJtg9bslkepb1+6z75g5hFZjlA3AunI0dVmccbutcvOVjoXtmo7No2kKv6eVEmyp6T8zr
dH8XJ6dEC7MAa6erdDVHfhTf1mh9pqQfS4+PkLJbzXMfOuTOAlAW5YqRsTj48WT4Y0waxJYYlcO2
jBcZZzpG54rirgxPdynQrTS8Go+Ga4njFlcVdlTBjoQtdv4ceMSC8EZc3vID6DGkrY5XZ9EEvv74
M0G5HWuUMpwhtshBU/vXzyC3/uTnAyYkjwCeKBHUDWNYtYXHRmUb5wkBg5ecAJdaiFuKsoJNFCEY
qnlGD9g+2p6g491MDqQZ+lqhg7IspQC99ICrc4kFJd8RCc82d3x1Cdw2d6RqAsLOUGcJ6UOEqmWP
9DM7mpZbofeCS1xngrd/u0twlF2nIs7wBPapnCYRnDVwUdleb5LYGYgaheZyyDYhg/krWCtcxofm
FgQ6eM1bDxc6YLTlJQ2+7kBqnydxKeEtitg8ykS3ntZLPk06kA0uclo4c/i7OLo8+yk528bqvuex
yGFNG8udBuLEvrx+7bnCLX032mhFiny/kLxnwn0ntT343ugKqIM3LccT5N33Ed/dyKveSA6teODB
OC1TVxdi1FV5/BBaxemC1oAdlD2yddoaMp5bjt0FKylES33oIoAuw7wQLWEqhA0X9UHBkYbar/1K
s7FxhF7pNZAQt5aR4lDitKcFIc8IpK351boqBkw5iSSsLr72YvLteyIhBdbi2nG2LNptlFojcjQm
mWGAF3bxboWJOdh2RcurUy9vZesTU48ASADGI9B/mUEj8fBa9rvpbk6Ts1MT8lsV0lqaESRWM3il
6+O4ZjUvv3zjN7SmQ9M3xoer4zyAw2fGL8+aea7/tS1WFRN/zhaFUh7xyu6Y20gWZyEyD6v0DnNH
Vq+wrn2qUYBeXiyb9fDf4hdh3waghfDKzfNJL5SCOgV7RAjmzDyVKEyylvoZwR41IzvlwMwpWN36
092K7lvFCt6NrEGC+34OYhdbO13ZSZD+I7a9m7hA5lD2b1CnNj5t0aUUjqStzILV48kXP0EQyqk6
+Db8ocE19D5j4mseZf4UZhPxy0MPDKWwmsAC19ipZFThGKZ1V1xlfdjhL0FDY4+oKUlxgo9b7HOD
k7E1qFlIjPBOcRALtTWxjT0vSSIvQtTf7tJloCHmDRIn8al7el5W+kKUBlcxMfECweso1OGrQtgR
brAt/x6Cy0/kj1WYAMUPb7fcx54ZN11UPcC2qmsKr8lBYw7/1q+dCZw2MpLO2cbVDkkc//mwg80a
KcPN/FdBejB1XdbGXS1U4XmFBiExUwJanrJl4wejSzc2eYYQ9SAHdFscWKHezP/o768Z6ptocppR
LpgFXw8HSDceupxJo8hfIlRzwGtVWWnCwrKqFGQnIOHlli+ZOdZSdKZfRe92fA+itLcy8Gw9VkjA
bfmhh8jjGMrAN84I+v996fsHiY87P4lq88YGzAK2H1aUj46w7oy2t9QqRZ5El8CrD6bfhbQI71Fp
CBXouptsPR9aXu/kzY2cJxyzS5svXXqQ09R2fcN4zMrkZbUGZq1gJ0nVYDhV+5qMO8BBnQiDHDeQ
iYPW8e7447T9Fc/69kL2JcV7XjJF/bgi5Tz12jPQvMWSk0fC3z/3Gs8/Vusp9j9mj0P1r8FvxWoH
u9kwCbR0TTOdyAOcDatby+hY3t772ip1Upb4GKyGVNa1ydWmRfYGUTHlothjfjPVnwnikS+J5wXy
r0JI9amH3vB9SUmY2sfmhADVD7q5U8ickG4kx8TPeIz7y9JfMu4zrhca5Oo6lgg3/aY+FR0W+ExI
z/GrwzjKKtsXk+QPCC7FThGd+aTBV6ePmKQe4K37MwssOqYmx3jB1Q4OxiSQwnJAcYypQaNfX3Ru
p1SjKTcWV7+gJ1dEo5JU9WVMZVk/OkZ1ccEKnKBzNy9xw2vdm3sMzfGZVd26KhGA+dQ5Q4PlneNY
KxV0gYYmZ7QUI9ll3plhkJD9mvsC6xF2HhqUG57lsApPshSoSy5Cq84oxQ6RLaYHCfRkag4JZxPR
6ekeGJ6JXrkfUwagMeQQDqr2kqXdGlEfQcN2Tdz4o2rb4NYq1ydvykVCtvke37nIeePPF0VnPJeE
6/PoZOY/jJquW4tExhqpb6S3+PczzklH9G1vzbnLxFd1r/WBMsOMZbC1DQM6eormQhDLh6H424ie
5Wb9a5KUbPmV2FnxlG7qvVkP7qTdf6C/P/XzhoZu+9Bm1OfYZgNfUIOvFLBjekSLA8icxpZ9NKyX
fFv3PFsa+1YXA3UVFrpZo7+br3uSLC9n9/tWI2TQzxHF9qpkgaftEaeqGDjPw0sMBBKdcjbsg4GC
8Yk4ADnJLTQIrknZD6uNuoXG8jfpAbyGBu9s6+aD9WJBPiBIbCm4WgYQOX4SoBCjjGx+nzBiHORs
a6EhlYlRKW1mpxbuoepe4WuCPKXaoE0NbOTKOQLRQP1FT0w1xKmkiv55CTwlb0ahnRVrt+v0gzRQ
h3kLoIYdeKfAjrpHFPpfbBwOhceKUhybXKfF3WPZ1Kz6nMkuOJ0v6NGSLw7CgA2lDCi0IRXSdsRA
B3RXaNRfukItJT+xh7Wb+8efs/y7EbQ6Z9jfkTx4CHO0iHJ4q9GzMzDeN8dqiNDAfvZCTZVTdD9n
H4ZJKfaZ9U16JhGMD1JI5V59pITL++RgJuNAeeHqG3rX/h2Duq9UCjPXMURe7VOLYrAEBRaXbx3+
FPP6rdjImK4ANc2BF4ld3UyEFMivBIpJYD4Bvqg2Id1ujFfd2j2T6npwxZ3jGaWoIelKEtfiUBDt
0JefWtaTje0u01rdXM4VQ6pXIe998BxFj56JDSEzzbXY4hAUPdlSIxFYtirA8J3sI+tOUIkdLJG/
bdQQSHHq2YIwAQmUqsc8cGjliCrQc6e8neT774/VMJQLTaoG6+89+wCrpqUhZWAB0sq4tTqCnRYK
3wkMPbXhymotVOKtWADpFW72saC7tLsNZTDHfwxXrWRSfvLE+Y11wj0h6A77Rcjq3AwV0jrduItJ
Dqi16zb4pt6L/7ksQ2XEEfV+kbsUFPdqMkBZQIQn4C2K2qXrxuEs4AoOPVRkBhuXbpqzvpicpF7+
ScaX7TalgzVOdR2OzeEqwNtKNujpPBxJmkAU3r5+QmYqLN1RYST/QSrz3WzrWUqINF18LnSfxvxT
3wJpiry76XQnhrwcpBteyH40JTHrbYv2U768t849HN5Ac2LcJxqYcsOP6pl/QyvR5K6GFGZtP7Uk
mHJdGd9lKDiJLkOjIJjlcatnQVJFZ1x0bjWj2JDv10EoNfrefcXcMlleKQgNw49JUNKezQv+1/S9
N9wiwANabbBsFD8mH9tdWzUV2uHmXvo4H4tlT5IblV1gD9SLwI/yfpcuunOjMo8aXmj0Y/qJQaMD
wNyUsn8feRww9I+6p7KIKfut75KcvFfDfQVkaWOZ4p1SSeJQC9xJVQETV3Og1FTWyXd7YjcrfFZ0
AkFThAvPFc1omt+OJe5DXY0fLnGqyIRnazyyeMTfEr0oscuwqmomkVit8UmozdJTS5oVXVitXdMH
c8XsbNPQL7BbGiHzCm9wC3PLjoLm0qno9dTuihLehAO16UQnOP4cq3cWO/8TnpiV0Ua2wmKQD0VI
c21gl//NjahXqTcLKjDbWsnnbfXF5zcSyiuuRY2wFzQaxiwPF2vf9VKDOGX5iGh7FAl4oHY5+PVW
TNXS82wiRyFzr+511PD0ukQGWbJG8+eikpdVZ5aY4EBY8a9K3LBKMBSw9CGB4aleh2IEl4d94awJ
6uGl0s+27x9koLstIJdYHVq/2TdQ+ugswnJ/sMLavK3WwFlznS25XVwahYoGraZ1sjlwKhXwloxT
wZDxtgxp00KJY0yoG1F5jfHK6u5x3Fwa/LGKKaGs14LGwnKNY8juX0nMPFXRNv3jXXajDWNyKe+V
eOYvTDdvJdfQzOlY8LVhN1hVJFww21uocTZfiC9xX6/6djuv/ixmAr5KQtj+EUit7ahITzEgt7cY
Oo02ZS5e7snLyVzpd/LZIMgOLY0Lvlxn/2Ss0I9e8bwCk9RLq3ozOqJm7227u0AgTvRv2UaNXdK/
+yWeuY1oPSe0sy/bAbMx4wDVPB40bUPcocXD47XQFvc25x2PWYVn3kNSuKhIMNM+OPl5oUxSB/Em
Yp6h4D4mmR08s678FzRZMdQSsesq3Swedk/e0IkqD22AihW1a5pzQGMl/WukgC3uwHaLWtLZxUHT
WpW47omDqnmJiIiJ3VSOXvUNzamWDdbO4olNS2FstDwf3717lmKGwcaHgRdIEVNB7BNHN0ktTBgA
WlTI9SVcmhMEkfOmUkf5G57+qzut+yb7NNLZa4rzFuMBl6T2wuKjMriNhp/9PYcrbuhjFe2lZVdT
JgUydv3CsxYRKJCz2iRbwslvyWjTWmnavJUDu4zK60Pamg/VWi2u/flUjDa8eBNPpac86SSwdruh
q8rxZzngxRkx+gm6htHCen29L6tGZgue8jSgl+HdwSYCwgFSaKPVRvnSqZX3FSOx/IBq9z3FvklN
6a+t4FrG6vsaEQQOzXmk1t8EcKof6XnubglzSHPH5S6V+6C8vOaHcjnVnTSwJSNEZtIUZTCkZ+uw
a/mbVq+XO/oqU0CUz3+KtcVKHBqyzGRqDahb85a9yG0RUTv6KQ0P6DKnFkpplAje6yDDmXri308s
DERiE+Tg+Ec07OcKJiY0+s808928Y0kdCkQqa0c0a62JVdYOzGiQlGgFnX4O/cYnwZXruEviSyYo
S4+5WNMST567CNQcVrWKvqLljwI4egDkzwXZmTU2l8C1ngpuBHbKwQt89s0SyAG8L9LebWeY28lV
Zj0wy41oG8Cj58M7XNRnhfg0WPR428lO+voEreptPU0HQFl2f/75GeL1gnSXnif39KTtnbl4g0nZ
f9UidVZ0JCk1rP/zI+meAdpETKxWt/Cx68KwrZ76MgE2zoZQn37r84GMJQbULLKUmXKT9kXbiIGG
TdhLZ+cgd0bQWjsD3SP8d5exjcS+wjTn6vRhq1DA2ZQeaKo3kcuNG/wo0nzd1yntE757jZcSIlU3
D4lOpOLJUPjj/JQsmfojadpEDjGk3g3luyRvE2UErVBxTMNpwiLQVnYfWTPpUZllztFyR24zdnt1
1wdGQWz4wMmCKZj2vHntOZm+2jLW9NV7Yo4+y64JeDBy/FCFvidYQvuF5QH1IXEXdmFGguqqWirS
VRuzDI5pULcbklDW70/XCk9YucvdQd3XnUVeFVd8CSI0F0LNso9+gKBhN7Z9jFwuO6ziqPqRMfAD
zcBJVMOxA2hvO+ZAVSZZpeN/6t96t+SFlLTz8xQ3UTl3bcQ7VPiFaPoDrrYzH9j1GkA1MEXRoJVf
PaIRdHoaqMbpF/2zHLlFRnQz89eNB51T/TTg2+Ikmt8rI/zlMgplQq1MlJxrJ/l7i0tCL45/Wx91
0VHbpTdbx2fcTXknk+IdEd5zAFpEEbLGX5ifLH5uy6fg/c9IqjY8CFcY6uK+fHvWd3qSPzzDak2v
LKrO+BKlBkppQoglmGhSae7743CAMpWqeCyCxWQQxgGqRekeUhF6kTMZhrHGukbTC0D6M46PO3+1
3IJf3eQqNZS+OR/yE1NqaQZOyGnl77seOu41+I9zjgl9I/5tSM4yBsvS/xZtzrAm24I8utFdUMz1
7l89ksmX2P3iUzgkVdFNUTmxAj5cSnStjVnVZBMHO8b+olbIIGt5T3cthal0f9IHZKTNoUjgKRgT
g/h3+tXT7ZkTSyltAyAZDHj+wRUP+H21ZDKDGZUYCJ2Z4KQKixjjIhJjt9c4Rao4HaJR7lhhvEzZ
OscNhFq1FGuDnuEh5TfURXQUUDnDsoX5/bhPxY12TErJeu0c3OwG6bSooGsggnDiBPx5hPHltEyL
kFU+pItuQD73RbRMbE+CH1etBNMQuIW7Wv0jkUJDg+uY57LMmXs+p8nXNQtblJ3zChJ5ECzCQqTM
E1kGgtfix0VGhC3sjGLvcKvAHsY7jKSep8IPhD2rnKXryFPEuIbYy+Y/vKDq89LqtUvf4sph/AQS
hb29lLfQ8Uo9heY0w3WLF4jO2ns0iWYFcP+R3KO7wo4OfvRqkwQ99XjTI+QKwWd2nwkVmNRE3jc9
250eztHRMZxQWL5roO8hTxkf0gUBUnPVFCzt33x8KC5xHrjGVh0KQ5E8VmHzs5Lwaxt783uLuN3o
x+LOv6CMaGZbdfjsVnlGenWi3oUn3Exyhfo4MVQzM2cbYK+37+fihFvncWXilwi1nTqVQsC00gfJ
0SLX//qCq/Ufvog8fRmNhBTMYMy5vwylw60lkqbhlidRfiPJIw28HFMptxlwxnM9wLDU8625dCKf
J9QRYHduHSMI0WzV9NdhtMAYW9Nz6nNG6XpIeQ4WV2i+4WJ5g6Lv9WGQeLkUoj/r9ut3Q8fhWv5R
M+BvdNvFzmT5MrKEgCU5uGlfwW+fQXMuNREIG/4Jw93Bp1IX4i6lOEgkEU77UPESoHZtgcu7QHJq
wE+njs+055g0OUE6MPCxJ0ei0RlwcTadxo2gBFCwfiVN8XVvptXqcfty9oBz2NGuDDygPqxadusl
N314PTUinqj8Qq0tmM0Phg99HrGXSOHb+Hd0vJZzsqpUW6OE8orUxdpuAYFzdBHVHpqKx8qTTW4w
/xhkzqhOhaLzxEKUvk46SCCjvnXXUA4IspOf90TcL6wgBn/8MAt+dqfoIybpZeI3yp2brukxd5JU
4g8v4bMxeDBbqAx1Uj0ajLu0V9xdktTGAfI9+9gWCuRN62gnvhkSj68z6xveE8rvQvrMg4LZeIn2
L0vU+uFWuidK6MDWCJSrcBgAqBZ0HLCTbE7YmRs2KTpt+yPBxhZxZQtyfj2AZp8ra3toLQS3E3qQ
pvOLufOKZhGppUCEKx3cuG57x4cstAlKke6ZUzjbbbx1RWcU/8KdnsDY2/rLMtClmDhS/XTHwc+N
1/zR7/bLigsyI3D8JnqJno7UMX48DRCiZ6vV+NIa7z91fBrHfvKJDPvE6oisDrM3OK76jzB5PJEc
NmAaqXLZXFppz/vSNLKtarzwq0ZB4pameNLjqjTqk0QQC24wbE0Yc+Rc+CiOGByzNhQWkJp8f2pm
ezWeeUaJ600CwIvNd+4/wNtLTct69kxXym5/uZvybP3I+bVe1q96zoWDREaC4L+n65ZoPdUo3Z3w
dwKZ8bQt/KWTcVR2aKZr8lJR4xfkDbVpnngy8uQnQy78y1uosDcqyjSrIpDm+KYG5wiLVkagRNtn
XUlJpQLI1/taHrMnNwvzTuVZLFCHaAge7zMcNVSH+eVBjUJat7TOmn8R2OMLwY05eAtJw6vzVmm8
GUIsp2K7kqcxeTwzCdrlYXcoVPn79PkOsNzCa65PTFoaAwB0Hy1zF6OpUoSCQodw+g4nvjJ3kY83
HhyiHveVLu0m6R19D4LyRehoiTs7wMVo7V+MYPH6i5nLfaijEUuVDqcu7nsGsbBgJPVBs3uKdAl0
1y/4c8rk5uWYJvW28euQsBGSjdXoU8dXWHz8aAg5Rp+ZtZLNyOwrmIBV03RY4iAcC0DYBlobobDF
sjoq5jhDGSepmq92oFJoG6brv/4v37JUPQ8WVsKXuUUV1hBWxt3HYTkDxNUVnz+sNzLtPeduW9vf
/3b4EE0cfPr4p8Sn9OvqP8G26o9i1ADdjwhR8ehfpilbAfmPLEmLkq30E3idrk0+QZkNN8FPZhHs
XWO9SWrpdpcLSgJfIVuAavPWWbrF7p0TXtjNDfk5cIVagdSHhz130yLKwkxZ9mN/VvuiSW+I4UpB
DXIon6enQlRf0xBo6ulwAqzdaLROHFXx8haNbGn3Aq7+1cD1N07Kpf0wRlsLBKNr1VxxZRvY8TIL
kLVcO7fCn0NPv0DlRQPhnZHAfoZ4Jt6XX/yPcxEuG5rarZfDXjW7h69KJpcoTPzdf3n9ki9XYND4
zHKgaPZ3FbpWjpj9UsIHCxiCDXfBp0IHUAMEPprNcTMubA/zePY5/YNc0cToNovOBVepE1Sbqm5H
jj2Q/z2RJQgiu+F5Nwxe61odfye5U1LRE0QlVzl4j63optnkF6LU/YYLu7ROmpszZyfpQIM4ChVH
uVp2r4b/O1i46WR5KoWuuDu1X1QFlaMuxahGFEUEMSepZh9Zqoo3rfWKbTBaSAhmhuyErMlflSBK
alnBJruLv2Cn+k0JNh+NRam3uem9o227sCaZelfZVI9s3kEL2dMGnhb8IOWZ/qTIs8GDZtCD/97w
ez2O3Js6JIZcadPfK6loiNLm2zAc3HX+r6DxubvL2GpaRErcGPxC31Q4rIF34MQBbdouLWclQZio
qlfHugHxx2rWxvlTZ7a+7pJ+8wxSUxH/WTzOa1SFabMt/9wx9OEfMPsjn16BlsiNkVI/hUBrLL9Y
u7nQinlJQVCPugxAFXDYZDWxRSQn2DspzgBLX6ed4AJxqPuoJBPAKEaPAZtZ3DCrWn2SRe/abysm
n2kFdNaKNH6HjqsKWPH5lwD49QGEsYNEr2ITLR65wFGmXYzhsVjxRQcec4AZIdcrgPVukklzxuKw
mJu917zy3FQskLTHb59XrHlhSJHje3F3dKkHh4EEvUCYQvemfS8rSU46GZnxHEIwiE5pf3U+E5RP
iyVPkgZ2HZC50VFHDfh4VLX4BBposV0OpNSRR32bWZw5iwyMKXF182b0kTlpHAQdgEb2DhB79+nn
lmCbsPBmqDwI5z71N99q8iAqLWDhH6CVzBI9sv4v6yi0R/j5aF3Px5uXPRi4U7/Di1AVg1PzdeC4
fxKbYe0pXBlSLcIbur36cqcJnMSJ+wB8Hurb48bZEZaq5+PmACvp8fZMjWVGuEFPrAP2pcvSL/Su
U6nDMzE+S5cNRo13XHoZ6t7l988F0VdqQ0wav5UirAun1fwjMqdgwxg6ZJiHGUtdPbSfGOFWDmq5
+RL8ECZwO+v4L5YjWG34i/ANcEZfBXX/nll01M1FzQ7vsXBdJYOR0QYPYydgLUu/8tC8aDA1PZ3G
A2r5wzGEOMSiy0c5gfEWbuh6SaadiDGn5LuAF56EXlex5q/RyhwqxqI0z+WuoFYlcwugeaTHDZJK
B83kZcz7cYooz0XIFNSgosrPgVZIATrkRGGKCu2fSks9muQw4oMJkpTnYOORioSn72XaAfy1dw1q
2bY3ZHWrB2OQ111h4rJJvJI1Aa58Ag9yPQ2BSnzLCxQMBjvK81z4XDWM/5gGvSVoMW2hakusELIz
yV+eLB2DYr+aAxoHyKvODdrkt0ZX/dBIK85lW/bXmB8+DE7cQDoFM3v5M7KovCceVfoOvTN/lQmf
YTi1BJVoeqUFzT2FZMqvCyZjyYo2oO3DsIqGWwl+4aShrsTLI1nhGWTQynBkZLMyQVcerCWxdyRH
DCF72dYKpO9kvp1dvKjEaICWYw4WfHxnP0V4qrFK0TW/1EH6pHaZ5o9/N0eA+1U2LIvUcnk9irfP
RjkXiBxoKCAbTaGXnGR2D4V4f5mPzSVJq7ggeuK7bwh2+Ai5GpP+hl13quqq80lbuiOcxZj/J812
Ag4/7KukCuj5NjNuhPPF1kCoXPHWz3GQxaAuW3bdPdvlsM+oG+Ju2w9S5PN976MFnbMcRSJflm85
KthwdoYYvObcnGrVvFyKCf5AZDVq6VALzwDd6zKQQ6oeXZ0aYJblE11UG0W0+HNTjtp0hc1GGG1p
331UcoLILlQ/OeIxxAramWw0y4VjsS1mb7msrpBU987XvAK/l75Lui+pMh50G+W4iJrAGI8PY2Wh
QDApW9wye+HvVqqdGNI/grpjp6P5Vqnb2LAJm+AKBhfPELnQSpVsiJJUT5wJoUK6sDJjW86WJQfc
ZEnhiGwdJcp2yq83OvZIKp4ISqBKryVBXLN9Gi0/Iu60xoN4xm5dKwitmK+hRAnSSAQUkS3QryVs
dEpxjdeA4wQeG7F3oI2hTUQ5OpNYcFBpPz6fR9JGdzA/h5w4RXqwal7jq2MhcJUUBy5eA9/4G14s
MDqv3Ofu4ql8w/KPQKUI7DM2V/zJqAn3BSVjb+W7aGgV1kTSixYlwyIlNowzSjFufRDHSkdMN7v9
a/B0dqdQHcxVWjfTF9NlRqylmZzKrRtzCwhymE0nZBz+d6TW5Iv0ZpfOw0n4OW77gZjOsTr233QI
fAzQSccgovJdyOTUnfo2QfLxZcn4yMnXZLv6EaLrdZkhoaOgu9aIFCcwVyah6R2V/xiKelJdLXwx
TygSzgLTfJX1E5adrir8AXoHxEEO5k1De0slwQk8csD2vzkAOfsT0kyY6i95ut/PYjVfti4D5rje
vMY9a2a+J7Mh5Xow8g/849/kQqNqdrVtcVDWBCJludruqEaO57cX9EuRkuqvilo463CMci4N73Sk
Ht7z9WsOruH9mi1o6+Cc9TzBNSXsjY+IMlKBKQZSHhkZmLQ4I53puwZqJm9571nkxkkGSOTBv28r
ip2N2bBQQciExfdy27miULNNOL48AhCKS1IgRhCutSENMIWKi/tD7sPUHxdYguC7hhe0G+/SU5wS
Vyp5qCIbZH9qxbCmk3TgQ5jGxEvgpBsfir+jpfyPf9/QUXi9o3Xr0vzA0A+43v6ZvQgSoOZWedGs
+VJYFjmDhNFOBM6spY6SIeiHOU+w5gPYizrrYFdbRVQClCArNNZotJ5ZO80m7nbtlIA4gCtRihXG
5xPOueUC+3fYU3oVfGIC+ZwTgEK6eaecr9aIA7K89C4TIaJ0k8TCbyc9RS+ygZsnnLHUBkDFAzBp
nWzEmquT9MU9OlnL15/160KAoa8+XRWGR/iiPAgjXmFtQPKi8Td3buKx2ZLsIbv6brDaG3l+Ml7s
eDShsuzQzdqUvuDnkKCE/NYIrrZ7RlbM/jT32nkoaaDFpoiWCQcQYlAvd9s6z3oBTP4+yH27JCma
+eeT53Of5IgJoyPbfxajZ3eZtdEqRqzbPpSTpd7DO82dZ24ntdyL9PU6dKDSUaGBkJz6w6SelR9p
uFEG1kAD+72573aGifH/8fAcAwZFmZsg8wR355R/H0cwSkySQIVVFp+xW7T79G+HAdQ5yLk/Y/n6
p88kz9EsdgYWo6U3z+2d9W6wEIJ5sBRPI2zakNw7aROdnYJ0lguxBRtaMq5nTk2/gJgKwaQJmRqc
ULv9REaDm2+IqLHmd6IEoW/8Sfl2+zyJAcO+S6xB92RFmZQJhtck00dO/0Lqr69nr1O+/gEP8S71
xnlAa92nbejBIL79PT4DKRaCXhMJzMwNAUvo7vm9AYVAmCkeYmpWLBVDDYFQ5zIHXo9CmgPz8ndd
YlE6f50gkS6C4xhh6P9uI9IIzf8SOEc6nzW+AoiyaKzzkkES/+4OznQh04aX7Z9zUbbxBItDTTro
u6r1E/g62yIuVieBwXR6eVnvgK4L3MIe7o74TWbktRcUAIYyRGpT3KgmQt85R15bIwoAnMs/nYVt
sR4R86VQoNALnYtuc5jqQRIxbtLWA3q5iFbSCuh9iZuzwLzG36bytAFrDpWmN8DJn0QpGGeI0tSE
VcSzQkt+mXFMZ7kMtEoNVgo/0Le7+vd9FKayS6VxE+m3aoFfMjkqbci8xo5vlt5cOHT63DJuH4cI
rxvAynvqbR6Qrc5Luv1CaqMq59T4oAVhH1s6pLnau4iWxb1HeP3mt4umcVJoAu9uJrx+VBtLw851
NWt7miWnh93Zv7I15JerNQmpT4dsHWIkMY4joJRYj9tcY30ejAL7i4tHRrFOKxIzKG5ex7NP8pL+
cn7Q6X8KyQZGzaX5khGsy/4oqUGyNZOgQlM5HeXWpmbw90AHUbFEugIQqD6k+3NLjclW0dchX30W
NESjRRoTBSPtH9JqjGrwR6mNuGopdB/fq4kMxsf+ZzD1rGkbTHdpPTSjOUWiFoFxbaPM7J96Vbcq
qQglGu9zfbBrjOZMsiIQ9eaTFvpOiyp2U1HBLil8mCk7231gYsXL8q3M+b8I3d9AA9Qjfl2RD6Ig
taWvTLsdtlbgmEJEaLNpW02tTT9UtjISMAKcocYMPPzKCKN/yRBeNiZ2K7OxuW9A9JkAaaxhACca
U8UdhXMS+5zyiaoQkKq2KDan0ZKYE5z8wM2pviRlKgMTsryNYqbSoMsxJYrdxglqJwj6eFBrGqL0
mOFydk/noKbNDROaH69L6sr/m0RoO1S0FxdP/YC5xT3ERfvu9uiwNi1JlS2rzj7MsYydXwg7Kp9K
xPMZL8+hk6NEM+N7ZaV5nLtfdTp0v7nyax1aLBjbkuTOMICDeZY2iOkcrkfIEKZjM0VtGM10w0Dr
nDcs80lSSLTeVRR+GoBG+OWxxnLXXT2OyoJNhwfs3xxz4ZXVLXX+VSWkkjejtj3uugGtyf5qZX/u
IvZIJ3NBhUBiS2+YJuvT8fBMGkZ69Lun4BS4WmE5rUiQEydSOjJ37yHBBVeGSqKIbf2EPJD6zrdQ
EPXG1RjDKIE59mzsNJpUWDlpnFeOWsMYEYqCzhfSEcSyXHNxu/s175TcywbXVlJ0Dhi+550zfxtx
4rNUc+NfZ8NLl8JJ7d3wfYQ5665dKL+y51YfIzhT/yb8i7crP8RB0S/rU+b5smK3tKYij6MIB5Ii
qivLRYX2y9oQGI9ibLe8eAujQ31c0AnT6id3dBaqjPX/tN1AsR2kTnrEhvAD2if/89bwNSLR7Vwd
dccwPbvurcXp2tDeV3YgS2aemxUt906kzQ9SPj/gdul/Cq2EYwWUrx0oJMrXItO2uRrWL2b78LBq
ovcUOXg1hfO5nWyjXN8hB5GabsRY5rCBb1a51x/tEi1XmUGJGSvmkiWuE4HcG10WyVISQPDqVmJD
XxgzxCXrf8eM/snSdUrCZPXlbEqtKPtJmGoAZd8t1w0fMbR/qj2STn30+XW6VttNZ5Vzf4CM22PJ
QhYww/y2LTl+QmsHjdQLMpPXS8z0k66/4YPKa3HkCl8WoHsjLufG5BY1zxse7Q/by0qbv+yGERCE
xJD59bY8vLRVIOSHTzXv/3L8sIEzRT4CBkM4uKvDV6yCSeOeJ9v9Tr6jsPLW1Y8Irkrclb7Th5Li
b5yizmsn6KvWjX+hLSLqvwhAb4pw0Sq7ckTQ8jm9dOP7ZcJeGN0XXyJCYrOm9A9GAOztdk8K4Qg9
bIkqKlb4Uubjgqwljwj1e6rk3QwV9bOqVguHeb26aN45vX9PiyjHzkRoGJvA0NNAF2cRltaqw55n
jeIsxxMc5jNwP/n0yXKFDn79ernoks1llbvdl1G7kzthpESMb6gURHs5cnZmM9nxfwLO3IOEE9fE
2YOb5ZZRAUvAXogJyWeGoYodcaD9wqVKUS390+939E6imNkNB3TfA6/OpvB6w1GGGnnBu8gP/53U
2cUXViZO5kQ+GCffPsZbB/lAsYCbrSw/FXKeef/OgU6iZeMqBUKPzHdj+SGI3fkALeHbdRFnLnkv
TfHaWdOiRo8cGLsKqOJoKtfx9n6r5RsB5VrwwYfp1bmhdTjjczZLAxF3JyYPw5KYucWjiVm6ch4k
nTw77YaZ1rqjHQ55WW6bebJIJxUdmCMDoWoUpVzggQLiqlU4kUw7/UScYi+mZQYLjOlRIRbjYNzU
DCPG0Z6gRwuASvWiK5OCqjtd9vgV+lFAH1wUxPsA40IPUqJGtyzQcK6aZ7IABGaOZp5XU3/9WZnh
7K1bUhNAq7i/lwpZhJjvrWsAn8pv1to2WLR0xXZoCogbUjizBsi5xZS9GVCRX+Fqgz5Q7q48eUiQ
lRkTjlosgCOr6AkvH9TIBCwt2nH37kjrJG7aS89mt5fBgZsJwwDDTK/4n2LuAm33Bbk+06H2eDGR
CpJ/OWRgT8LOwTufXfEreQ76UPIV92BXiHvYNe+kNP9CWFzqgTWHjmEsSMfvffPUr2fJemxBj9iM
YxNLWsPeDGsLRGyU7/q+rG5DBKqriiNQfG1XpjtJf8iJpGi47C9/r5JccG3H7Ml+JTbKV7M0QjLF
3nHpRUyTpZwQAkGcaZMTqtxcJAdG9oCa5KzPIth2LFSvB3BIbOF3SJC4uW9Aq3RAmErv/MWTrn6F
8kyE778gN+lUBvRHJfV9RBX4IG+fe2HKv7QIl0rhLQj0co0obdUbd1xclNLK75OHrmRJmvjREHL5
h77Nz7xk5ifyU0NxQMgLnjgkNFNTUqWtlfj1D7cRiyrWamxaQ+aqb2YunuvG6i7NguToad0MTIwi
BVOGN3GPWL5T30CNsn1swAya5SKJZUgGW7+IQQWhVzHxssEnDd5WG+XSe4cIlcDIBp+w3Nb1hj4w
oN59qqrX1zcI/cGALtb+Lox/lAjZMK59FTod2kR6yNZZhxBWibFsBymXt8PWAOP87Ac1tVUuEHT/
PsXhwXAbuFX7EtX0hn9uDJFuZe87ii+J+QinRHxLZZVYbaDwaZW0wVOqrMlj/5cNDtJhs1urgzKz
jl21sLP/bQP3b6QjojbrzhlbMEnKUZzpmVCq9dsx04CM/jlTew8lLVtC3gE5Sh6v9lELmIzqZgkG
RthxbKK5tpURzt4B2WKiS7h7DXToy+R3UwtuB9Sw3jBP1XFIwuNy6jl3Dr2FepbXPYRyyQ17uR7q
JTZSXP5ST1OH4UMUORR9zIhPyZImB38pGPOJO3NQvygE2FwC3QiUKIXoJSIIPs8yFRd0QU+DhwJR
3yfGgtqIALvmM8F5w1k21Y4LidK5LCQwDl7RosAIe5e7NATXiyjDO2y88sGO1U9NgNM69k4mN7VW
ZmJi+dT2sLoKayvzPkeI+EjP0/q9oWy96RIX3LVLwrQxe4khbbAQDwzc+8ZQ3oRMXrxFylQ0rgZH
npTwXdj/7pCFfr5AY+BGkkSu3GC34TLPGGtmGjDzljMj24K/m8ByM5Mr5gGguyDPsiqk1WCmA9GE
wRkZIUB7A8Da1F4HSlngQ6vbA8Ri+b7GxtwWAeHfnopOOb4DGeWeZWAzHFivfuvbou/egI6YHvXi
Bx5P3Ohncbx+H0CzOGEAvLnX0UEIg1QJSzIEnzvpB7yeM/7dKoh95qbP4sv/4nQboFMq9kdFb0Ya
cB8z0wC79tygVaAIzn9NKFEb3LAABEpawTkEWsUbbM4LoJ2fSrEECX45aQMRDsjZy35s+KYH4yfZ
fsRk0Kp9fFkkSOSujEPTsVVwkxrgkYivq5kXIRan90KsZWzfJG9nlcWCQhYv/GjmFWYFoIcPqYqO
LcX8OxsXJSV5GdpG+stT1LOjHkqM074WogweLc6fs7MBHkjUY22Q11asxSoXgrkw1bRgoSSlaVJJ
D11MybVlsMiSKgpdGS1OhSp2zCnxDVHWFmbe09rzH19KppdO2zAtHxY93q6BmLoDf0rB1yM4iqjj
BzGfzZVaNudsBIZ6OvCi4pALG7pIoW2o8gdjD6Cu0ORbw0IZA9/6t81Zgn2OS62MR1SMGOWm5ixK
GZRam8bB4rVkom3xnEmIC0rVLndtvc/ZOOCwDdzbb3v4kpW3pkYfJODyHGIVItTzfI6P8ZQyLQG/
PWExTqi/EAvwvPCUPNtdh46ik9xEBm9o+RGwTkJ/wXB4iE9wwc/5vs6xxG+Tb9SSK+06VGGiJ6Hu
ephTOH5bh1TN7Apm4KIREH3Pu5Lse86Y5U3hJP7ULOqRHoY1k/7AkHSv2pgCR/Mqqp6COXTxuj74
sJAbR4lLzCMJXhhspqBGKzHPsrnhUDCKW41LUfqzTKm7qDDv8ay5GfduPyPLK2RsLc60XA9/P/IF
ltBp+7344snh/EQZzGh/yGry69m/BC7WYTnI/9wXp9tOAQ/atMqmrL79aTCQ9kSABakf9i3XIBva
jbd5nkAKp7zKlWmENP2YPyqHo7kpTKu12DLaxuHxLB5Yh4dxiqn/cpL6OoLDMbAffRgznQtx/0q8
IQmEXTehBD3RdIKpofTNSfXVBgo03ePGG5iOUlxkzY4ur9gCNbHRN/SHzjx0woow0U8Cjc2P9f4A
QGOnn+UF/Kaw8t1696gaHMqdtot3V2ss8FplQ5OanId7KYH2/Drm8jYr+2ccUIT19AJNGGMVm176
ApjkmvBVTBUAqgC6F4XoZk5WNOd+4/zrPrBGBAP96s70ZshuSAxmObqQXgDSJhX4D3qTKwLdNZ8r
p3gvsq6OL4DnSOUWo0JPWor7P69xbUKsK3B4fK4SPkhH14J75IaWsFtmePuyCVSKM8wm0IwOgJCd
YSj8D23JVlaUBKqE6xAHzIxHXoeo6Ub5Lz1pivBCPbZ5tHu9s5qOaq/NUSyNYwAaDbkSyuY2/G1J
QdLSiTeV26smjygY4/5i3diEpFGk9XMl+fXOhbAMP+a1E60US3LFZFJ+zsoXlihhibVpenr/vQM3
d23twMlpOuLKK/jb+CsghskVuqtI/sMB50bEuHB6FNZ/usCVRrjgiB9QETfCmgvXNdLV61rRRApW
WVlsVhpwtT6yrFKDlKShm8bamljAgw8lvj7pi+TV9kzGlqXMH/zNCW5XSfEA3/FcCM9t3UsijECo
3R2GIDkvpFINqBfqdJ6QpzvruxA6sRVUtfEgCzs9N64IKSXzBk5yX1FkqZNY68qCQEfJLIEYq08a
+kkWrSfViAqJNAPN8hidd4zOmZSHqSOnRXlP52bxLbBpVVaWNgZzAITz7C0prNu5EbQ2v6roKDRO
ImtrtQXiICAm84gH87Wmon9EFF802dVqQZWc54JtcXMe6XySJXP9PyzL3BR8irEbpO17Dy8NbIJJ
GXH9ZtcVgH99bliR8SxxDz/ukpgKTr6xY1DZU0dYAw3ZGHkx1QcwwZlc8zkI2eVfop2sHZXbUNk4
c/w6i/coZyfwQzVBqn/6HurqywaekvL5W0N5EsFtkeMBZjv1dsdo74f7Ec9j6bzEl/zwc4AiVTnr
XfzphukAShPhdp+SkU4Jz6MSZm6RjVv7IarASITlZifGgKkI7b07S8J3XHwQ0nClnO/zLIKVLKOI
oW8QJxyU58xJB1AEal27rPQHOp3ylSg1Ry794uoDkayhXOK2I0CrdGEYP/HoZPSc6mWfE+YwvMwn
UblgzxMKRp7J5sTWNvXwa7c61eL7qMogrK5RoHz/KXQXgXpYM41Xg8UrsigSMzTzsI3afBAHrMew
GcaiaBIsLPvpxGEKleXjx/hROVQ/1B/6jjHWUhrtsRR6V89eDEhfC00a/0xwrvLTJnxJLEDmxfUm
GTAI0nM+eN05QJbBS5kdP+fm5KkDisw29Cu865IVX/d10n3apTLoBTbH4p80UKbqHt+skdbvcEYT
rfbBzSH+spNRljbm3ReD1EeKPhyh7tE6itnR903QAVMrKWtxsiCidnXFQezRHHtcKIPt+eqV3/lJ
GF0gYMUevtTeaVUmH4XPFP3aKCOG3FpPr0ylIczWtgTfq4g1gdo5zU6vKN0Vj6Eb8ifGMRSi2Fyb
moTmJLfLa+y0KxLu7ggqBzMkIzOHC0Hg8fWyQDE+0LXxB39EKk+8WqckT6r8Y62/tdk4LzYrsirz
QnjcKEppnrhHaIhZqpPz8vcpi8sDoiqJZzXv402WQ6XZ0rHvoTr5m2KU65gVvkOHsOWhuDlWsNMe
fUGNHnaTCO588qNuDP2IVL2AlCf80y1OXvRUjEDtW5BTzeQfMLdVNRsINMuMPf0C9tZEX10Lz02V
zxn72/2LOraT5Woalin0mi/B+byu+E89BHzBAu4ro3XXm8OhsC+RRr0wWSwoaLiK3BzKWtNsJfN5
mpVAuAzvxD0Axb6lt9kpy5uD7puuh7x4LFhKiFcAwAOduuh6nFrLxjjskqeYKc6rxZdWCNshIpF1
loRnw+gZ+aj/h4Kxj9saVE4/9hjsfXA2UjE995mKeSdm/N92M9h/CIqHh4D1T4WqTKVFEMj1n33H
ZwGIHVXJaTHBe6XmusmyKd6ofd9sUpmJmap+3ia/1bad5uf3VfQohgwaFUs70w37kR61w2F6PPM5
plG79LeG+OVgxMD6CGrKGVh3+jPRulEMDs6Os5/nGj73gblqqnDpyWXX60YAU8lIfkwgphqid9w9
HK07BbsRrIJGx+mJy/fGpnTyv3cL+9jG/XdLC3uPUnl99n/aSAPtAjf+YAGIgQwLzvsnfZnXtQpJ
hkl6G0nAu2By+lYvcCq09CQVdVAcwOyAiU9UqFDVBwy7aKbHIJqOJZcJ5FJipj7mFsBT4y4lSfc0
81zd0xFkLBzzXRjA9whmC9k1/nZvZIp/fBfCmHEH7CtlO9FlMgw2I4EjxkxSkQHPA45rzLsewqIc
kgCgKXeTsQ069vaK2uT19ugphYize/THtRYz2w39TX68OwF09yKXv9FShRIyyFdZha8NQNWKu5l+
1CDQXja4szXS3OxP7qP7KdDp/siPulyxGFWNJtFn9pzZ5cy84N0lLowY3+Z8/HHsUuOuGHWtu9dr
fIceLRUpg8+zgok1Wn+ewxz4EdhhcnzMaYEkfrDZV4BJGk8tNHoUh3/A1LVOEJM4ZgPGRKLbMoPD
1WZ6qufC7Hl8ieIxe/bhko35u0E5iafobe9p7Kl40d1xHhhzo5GR8M6+nzsLJgk6uH0MmPcfzydd
8FtC2+FkVoAmO3yDpK6IB/s4KHsixILpy5meb1YcCwyLAs52xItAGNONvhmvNteLmCnZuI2ruu5H
ipdBV2MANvZTu5aqOQCECxLh1n1m0lntUMjmagRFiOUWCai9CcUiABhrEyBE9jy2+u1pcztGGdTP
PJUSSEqGju+3KtoyIAxldqFmKK4FPC4eLtc+GqwPyNK0Kdrk5ObwBxHNk5jZMN33+Vx1yUHHdgp7
1z7S6xt6Vkpl+xccRYh+ckp2HH/GP3EkBKZ+F4L2EQN90sIxGqx/5kz8aGh+Jellsn4XQvL2J8KZ
OM+5FO42dwcUTjIMM2W+zh32TVM0lkCAB2sN4ZtHcE/dsa6OxopspbP9opRqWvPtDy4BIWf862wu
ndyhfz/EW4+OIgqSMMkxwat0ZXQwjtCExKgdgxWbzOUyQwRtZUbueVRtyUyA3+rWoHW7CPmYS0xo
bV2KB4gT32Bgqzmc/MoqpklYLDBFjfucXFF0UnRa2Sgu3+PrZ+N+8IxYxnf3qQa0+xple5GKx8CK
4WaBBrVVy6eNCRuhQXmx2m7mjGU05RSzKfqeom/edjaUViZuOSXKaXlV8db1AqgIrAQQyx1jS69A
fTAkMTNZ5kqV1Q3fGwLEd5Fm0Uy+4VPs5EPj7uhCn0/rNVgS6jOAhwx1ff5TT+W+rh7sI5D2ZrVr
gZbf0yc6Rk8Bu2EkUUhussvxhxmF2NJBxZgyKKFrmLlJi1wlgttTIx1Uig6b2Gys3br79b2xmUtV
KBBxdBFQeMvgi1kJdTXUjby/LH7kGZ3S4ObCgiZvuxOBfsqhEKJB/112CFfs/WPJqoONrdSa54Ol
m69ml1SCY//CL1Xufh62REZaT22QSE0dAdeMFInDjQujmvDabyP4uy4KU9JEiSo8zT2Jez6LGk/x
tgXT58PPdj7vaBzskPgYf493SlKSwEQm3JHOKrxF/HcFTfmnTlVnNAai/B5AiTtHImcyC014SWi5
vGjo+rfNP89ttJtmzjEYABtO0K1fk0MaWUGxYWzEOx5siv6Eo67Vye7CknQUvnjPhZ9E58jsrjTl
U3BrN0ycQlT2jYCk/snneWcyCE97lfFrm3HVYm1yzCeV4V85fcufoXKTm4vD7AK7HUs5WUSFNa99
fkHVoLVCs6T9TRLtkaZ95XPrz1eBMG4Fa3IQrrnuyk5ZDyFx2c/0QOZUCOVXTIHFUK2/6vaQVORT
014PmFnl+PfB/kMaADCgUIwg+wM/jtRrSVariDGEsXoYURkx++CpC6Ju7lZCmjFDonJE0xRTE66u
0kFdEXTZN14tYpdKvxGZXdMHOlvItTlg+1j4YBAGwj1bvnfT6nc3VrO/ZcbcCbdQP6OuiFx0xZH7
Q5N800gQGl6PC7cGinS745bAi3iYJ5byY1Ut5ZkT45cSsz8kXV9Y1R27EvQ2QgzRyR3ls7Qg7PKq
EHLGgflsnc+rGfp1moKb63D42BapPhXNq6WsiV77Cc7leJihRYo0TQSY+mKfnvwSZGaxe+EEACrn
8+7gPKyRXg54iLNm3Hgsq/AFPdocZS09d54QlH//+nxtNpBy1j6dRxj49QNj9D1VLl1BYWh+EjJu
xvibE5rRe8WHmoLVglA3jLSInY2hrzTtmZhzQp03funeTRWghCnmdcgETdU54oQ/zXNQdR4Icn+x
aEFFYmmnqXoFYkMHFcCDy0mOqSNfH2bQZDWstZedUlx4mSLGK2OXIkiSW02M5EyigFQv3PqcqSmp
UE3BqLOKO2QlSTdZ6DVj6METhxFrEn/D8VNoMNGxtBKqTKkmRMxVj3jnu2nHEFX3be1CFwPqx6oZ
Io5K4OuR1iVc+9H/D1c5BvUPrBt/deOshTpl52vowwWqKmE2dbEWA0XsuF+Ks2HiZSxP6GBwpdtt
I1axRScWr7C2dXx7FABHxOt2qUELGKNkccSgBfcqlx3F9QipHKdMViovA7YvojNDOD+uyLVxKIqq
6r+1PbAhJkkayC7BcenjSXNUEM9fVmcEiXujlbs8zeOGw1VTlLccKOApoNBR+goTKb5xR9kpDbIZ
1HF/eeXFPT8KTNJ3UumjL+LL1tAqHnrOEF58O9PpVtYEO+kDDJtMmaCpTNWzDmhVIETnu036fbHy
AxQzuaWkBGGpGQIesJSByzsP0Djf1w5yBIvyTo9gcs1tWCMCM5UcUAw4jsCpTd9MwDIkxbCp//5j
SaAwVG+zqpzh5ik1R739Fn03XyGLz3WcUDc7C6HAy531ISKa+BsYY58UhWRat02dtsbOUSF3Z0l3
jo/TC54/TS1xa8P02QieaBhGF5rHaKv9EPZHF2ll/Rn3FDtNTN3k4vNWjv25GNv3rOiS2UpmlhlC
SdDaV7o5/T1eQBEMUSyLSzNeUFzar6mFohUV/EdgpHhvc/hZ5fEtYVSbnFHyZqQTthbnYXcnRhPw
+kNXAl0EvEV071qdCizYyMBZkCyQFefylpmrMldztz/thGKiEKGh1d05T/pa+Ynvd7BKu6crN60r
lZRxrgPvwxRnp9EwEHE4aBe+mG/OA2tV8tpfli1ygBnOU3nGaPlc5+0ERHvEIryDk9SwXfOE5J+j
TY+s7ATaa86vbn125P6C+kQvNBeGtuxEJ5npfXHoHiDP7Ltug6jfn+bnPi3ng2nazlq9cWDhe0Ak
+rOpReF0RVdkS4/Ub2pnic534frIQQH4LBoTJOelT6QsD5BwDjJVE/PQ8aQy4KI5lBvMumcvRYM2
4KShhwrcJ8ov+cDCaJvk80KdASR3/RS3fnPaiAm8SHHrlxeRvrEZgYVkvhElUDqhL6nWaa+o9dvG
N6MRx8TVqg/gPVxbqnoIRlwOcipuobf7h0vUJHrvzORxz1ziegjGOPMNF63WSb5qRIPprwcCZhP3
5ZvR4mSByw8WTJTSIYxDy4/kUTvuJDLMtelkBic3LcR3trHBzsSwazErau4NM3beY14rjifrHxyK
NPYv+pgle3DqwFUAjzqisUTjVQ0pQk/rjAKtnPjHewaY0/NDz3wJqgf23y1ADaOTfWvGtMLtEFHn
9c2aX/fS+F5383J4KFUtTORGQ9ZnP/PNJIuj85a1SxBFTfDmAi3B6HTItnpoyz577LV6N3ZqhFup
T7q3+4xsYLGshGTxP4ap9REzcUXW/OpVxHqScwNea07Kgbr8wNQzaCPWlidtLi+4UwG04VXTY+RQ
xR574P9KUNlXZcp2DbSRn+M0rOpOw98eoJjZn4Gc9IqlMDSNjqVO/YwuitaUNcyO0ESiOUYvzfLU
S8+ErgGEOR8ZLBG1ixHxrjEgieXvtHK/Pp0zXqjKfYQmXXvQtg/DfK0kj70Bf9fskS1gHkTVLPYk
qtn+Dolp7jznzf6ieoiTtAsQGmG55epxq0+rb0MX5ksbSSYOhAmtaRnyl+eGnu0JW7heYs52KeA5
v1Q1p8yp561ScHLVUSd7Sod0zk89XXWTFSimrw1M69j96BbGwLEnSSnG0dh18mdGhhDLxBW9eqFi
X/KDi5j4SgYNAgH+xw8aXc08UNQHZRsaH9IEBU5xte4Jx7GhFkzIRMzT8XozssPLj8OGgky+/fwM
AYd85naJimpWFBTjZL5sd/LCu48LVU0+DgvmpeSpCFR8LGTSt/PyAN7dGv7i4tJnX9Yzk71OMyFK
mkfgHE4QIFCTGsK1MdzGxBqwlXQbEjIKr5cSdnwBziSd5H2CL7bvYIzLQIY+4rkfoeCJGqtxXYjf
4di6HBjnyZR2UjNoLHEvUCqlz+rcC9mDGXxcdffJHr2NOyCiJSAl7gfu1uYWUHOYeSc6zPZ1KVgj
r+krJ8h7JPHq+1rYPny+9RWbET1Mkx0V/rVTLf79FteIA5brGnJMiBlrLuWV7xzBEDzidufP1QOP
bQwiKp59GLLs8Dm4zKLHLhjsL4i69SKTnu39MUOI7igCsQ+hO4b7AFIK257MHTCFwBTbyZl3zkcg
UVB+nq+zJyfdQeTwsnPr/hHcjeeCleypx0OsUHFM9Gtd9Eb6zsmHxR79cuVEaWFAGIsnoyBHFHZY
14W2XMj66ra06I0aT30yeZ8JC3U6NnS3xn5LePkJ8DYwpcCRfDuDvB7kG+J1bqysXIk9OsuYQUob
4IyzfLwZduu8+4/zov/SUTqtxOptJOEhRv3VWu9kcf3eNkyYSbLgUz5jtxuiFhDS6mfAkpfiwceM
bYfSHkMrccFr8ZGhGp4/u3w7ste+YkTvMKGNy4VIih30ow3EOYWuRtSt6wYji1JQU/jSV/dc06Sy
9Rs1S7aZAiNOrWojAVM6lGHWOiNzKfDRm725eukt8TCE9S/rWfyxtEpll1n4+g6ROLf2J2hh32h8
JVh2oDLCqVKWXsIi87vxeCAToHsJkW5tmMmUd7grbXS1wBP6XvbF9Vnk6Kg9TG0pe85jGXvDhGOl
aSC/6fG66y8k8UmTwdKok2jIkw98Qbol4sYBEkUfcK2RlOxtjlVhX1xiw0jXAscvfdCdcqRCTDtX
venJOjBdB55PTtcoPGXapwPJfGfX/wUL0HcT7tbSQi/yViv/c/0lgeau64K8VPLzamTn59nBIKRX
Gx+jvZ6BTYuokY09eJtsSpaVqT2RQWnftg5coqzG8rIKWI/3dWcdRJh9qnzNQ7fgCR80hVrap/Hl
GDBZuSZlG6EHoRbJbNbQg0+F8lzlrJQzL3YpqmrXkUCIbdqbSBUbWGg+9Z8aYk2O+F0XlH8Hvsp6
kp0SqSeN6B4Zy2CxGYf8gWuI3TZ6u0v0O7x8h2jkWmr7CKMjH7860PfGrtzHNby/q+WaseP8t0iM
4/F5ANqoGQXnYKaJm+uwN69tXXZecsHc0xLh3zxuzIMi1/qUiTj61oCYTnt16DzjJTo8ZwVok6Ap
wxnf8/92KjyiWaiCl7Z3lJSjxu/hssih+zZKrlCcFk9kPxKTIL7CVkdovAo8oI63oVGKhMeZTyCN
Eu3pafwLTZZgsAUe5Q/rIcBe8LC/bIC4otM8kQ8Vgj67uE0rfNe+k2m6SiNfuLfORKFPFxTizggj
Cq1g2u0onxO7GXeuqtRYGLMfl5eVd01EAhVD9Pt+5TTnIxryApETk5j20T2RygLcUV3eFO7pQHkD
cf/7NR+b3mbiTRyJj7mZQlPIAkbrB2/UJ35IPwpjXMxRnTCiFXHiYhgZsUh8T85k8Ew5km0ZEHVP
LwMGwXx7Sh2QCPaedEG3VEeMF9vJddeLtlDyAHL92aYeqXp3VjW6k4ZbiIN+FPHyRw4A5sj8D/rc
7UQFiEMDmoutE1xpuwWiwd3+18zIprJ9iihbXPSI6Yyae5G/P4yCmEKBfjzhnrnG9F7hY4Gqf7rZ
P9qpFq6+7MVigw8+Iz92zN9wIhpemhHShKESVfU60BP9PScCqTIkXK3bHiAcANhvZC3pre3eJHy5
eUqAi1z4PQqD7vbSqa2C6UN8LWKZ/r3Tk0w9KfY7ieNmGYzNwCW3DxYsi3tPVexB27k1zy9X9pF8
LBHBu+HLpkJEoRimJ8Ebx0t82e+uzJ1afh8kcEyJNuQ+I6l4S7UCpXmt64AregviT2Zfj1h2fI3a
3uP5N/oFAYmZtDfyRCaEbK0lyGgFNYfAijllV9ZZj+IATL/dXAGbNgtmjlhkh98qprddNNxGwzlt
J8C1ftznMwZjOS2hYIqMdrmV9ucXBrr8L2g2gquBZq4BJAnvEue6oagQiVz9O57R8WlpVik3aVzv
MUtsof82TXmQqdbcJ7h1d2V5SxZkByVJY/ViV154BR6x2ShTDoLxBySEVREMl8UCz6s3MEWYEX46
l1JZ7pZqVf4aRceXUFi2xFuYca9Rf8exFoszkBTqjuo/5QnSNzrlpWtUyOp9izD9bpshJkqO+yFT
BiIc0ilCoNSDa3FtYClugxS1ZL56ZOoNeo0jSMln0eyciin/tqrs4Oyrw63CQ3uPvw9RTWyxogzZ
dIFu/n6VMNXPRYrdt++aRq8dXbFN3SCyJKYvkeinNPEWA/QSvi+IMwkleM6QFDbUCsvvE3BKIdey
FbzLd4vDRGJdu9n6itG29BCiDUNMo6JDq1S332g3U07DGT5+U0XxuA1F6AUSdCqTudeQmdBWW0cQ
Lg8ssbdFFy1MQT2QyC9gFGr907Rmg7w1RVwe3T52zC9LXXhBj6cdhgDN4wT1IxGMkR0ye8LJHpGk
TE8IKOoy0Gl84N+Le95tmeQ7GsWV0nLavuLDRif9vS9Fv13cy/lhfeQwqRNL7szFcxqgdIsr9qHC
dQDSylmzpFOajImJpTH7xeEubq+3z08oJnuNTXYK/ETOPcPObQjQ62Dnv7CKTTRW9mpSt2QltQ8N
VJJ6T+D0VS2Fr4GYhrffrK3f8rzt1dNFe9IVhijL9zQMokRpDbjfM+FBIY1qUaA3d+6VlF/d3Lu4
Tq+aLda+je8LmXLWSPyq0o8Y2VdtrF8qPQyV0O99J827nc3lMvxo9gFZxrI8885FNiNPF94kKztI
t0UuDAeZrhAICDtNhwRq7jXfXLE2SQAvQdheTp5e6ZJlVnaWGXCP4s/dsnzdyQ2QtkM59kNxsnDc
zrVGzqaVw8QY+2Jd7OvpLY0gE7SjhbML4wQeQmWPIy3ALg8Wz1aAX33EuyIVfOXPnkZGKR74NVuq
RjNSXcKui4vW0EdgKQ7nK9aaVB91uj1VPd+x+G0CEEsSUuLVumE678apzj3fU8/VBoWq4ACFiMU/
J0VRw++uRrXmRpmSHBEJgQaCjPeYhZBLp1xd6yEa8EunCwut7RUghxbKI7vybGwIBJ1/pjf8T15A
MSER62K0PksCSmht+yniuMhT4yQycJ/j/FdlYJ4rYkFYeoli68wMuSV0+okhw8D6hyhQ806WrErL
O9s70HRPnRVufLGHp3bC4yYq9Amc4VKkgn1eDl6DlzMEw/1cd7zB63yN88mLdyDnWXESPTFU6xmk
wQDIFGckm+9/K2RtgLwIxLOY+dsfAeO7PzG3Yb13pthYJlmZAAXSGpD1104eQDjYUa6KYGNXJYGb
vEh42cgKfVK3B+pvZKMwOmy16dkCbXP6H64R9Wu3rCoYTK/IWqmfTZuZla10Yde5aDTqGrhoO31L
w2iU52Jo8YzSEsTnvww5QJiREJQG7sn/KjKJ6ayQrBaB0/EfKKtsAqode/yzMTLzeYTS7QRCHfV1
KJe2zs3QTYTC0j/NzOgJDnA9MijdSgKaV37cR6wfP8GHtYfVkxB8FBTbDJlw2L4C6J+LxmC2iDic
+fH/v2s939aU8JemS4bVVVw6pv7tIGiP6AXFvhiWLvubbu3Nv67DJQXU/mvSTHyKVXOcRM9WW3WO
mFNs7MGvtoNHiM5gNMyOQ41p09XT9SlXwSzRaL4lQU8NFGhiRNDyzKNzo2KJZiHCY/xnqRLbHwRn
roW8C6oO3aI7SuWsaJ1uvC4XwxcLQR97sWfjauDL0ffXUMLb9iFd66Lq3efrEhtCFeSgIobLI9E5
XS+Ucgo7bpnZxrw5J7xpgkoIEHN5BS/Ys/v9/sjZmIymSC0KPyj2idbIlp2ZO4AS1yr332Nziv0d
SwfBe4tqRBjyVOAfbtijHHhXHKmbsYPUwxprlpy1fiDEEYcPYed07Np6X8fEOq5DkdpoX9TVurg/
GTVJh0DEGWlHpJGoVOX7gxmDScxioLCgBVu+R5vX4gNZ9zjfLblmQ2bkEs4AZkmERA7gOAv4oGxY
GW+ugRRdUoqLSiPb/voVU5aFe8sCXZ/KloR2ec8zLdpbrBwNd62Cs6b0H0dBm9NIFVSLcW1sZMWW
ucFV0C3+WQWE1zSa6VH3WKB9t4wnBcs31b1vYVGuZvTeiVqfZ5SR9WDsISLJdOu/1PtOtoXENdJz
tYFP0HwJUgLi1AseFjKreYUeCNJP7eSjoFa4ZAJSZojKDijtxBDar1mYQyd6h/Q+tcdvCCLkrIzK
d5S7znAJqLnvVrkeJKuagBXEb6XKOz6q2J0ovdTpryBEAnapGL7JViCBYO+nyHj+g6JpN71hzYTp
XRM3PuHGMM/j6k29e4BbCzMd8Y8YGPZdgHnlzOx7azh/x2Ar1eMwM8pVYcn+/nch3epJZrP9YU8U
JuKkgjn8mJkXbIeEECr1KsF7opl5QVpQq/g7jVx1b+rlj+XkfM+PxZojlEv3sLi3wXWD40JZq0RR
Gpxdug27+0Jx01ri0rW+7IPaYtxmbiwHkup3Yue2NSX5cTCuC/oQToC4ecvl7hBcwRCANuEex+Lj
wKOlo0W/IGPDT63LSKYDPeG9iylOp2Qj5CDDwC8JNL5VLoOeqmVIvWbYz/+FxIzCHTRcqKTvHvyP
NLiAJZ9uuCDm+YNGRDG73/WDiRKiRhxfKelaBkDeFtLzvtsiCQyg3lOYzGtgmUuezxXUSh1TCOqG
irypCZuZsJITgDMudXxhhNt5bLdVXpzFFD7adSsTGjr/6dDQ8+h3XsbxStPs0y0D/zOwiJ4GU3vr
TYnk3GKXpjQWxzRNOFawn/EeOYVDNk6VeRspUYMgnZ2SZoGD4ZT+RmHygsfry/WETYOpbClBu+aM
hHNfwE5wAPyxIE2bp39nrb/UtZyARgFjjoVAv/T/ORrnb2bg//XQ4UbN6xFHXXM4brW3DSw5UUM5
yrTRhVbzb6HW4BhDTNqVbocWOkO7ivcgE2obR1rO3bDJClS/TKzH8ZLqO3lwvs4ircyuyHsUYuhD
WrR/f+lP59OSbM6EUWt+8Ou5RwYNBl4r44VZ5u2sSoMMnSvcGE+axPYucfcEvUqAcM7wi+/Fl84t
AOIBqYW1e96ppSSilkpc+1teujRVvpftxsTHdO1l0k3Uq9lYLQy+gO4UiQPnsdng+3yPGswkXRQx
i0uFxGKVnp8utanDc/FY0zyLd511ZduzGm3wLC32M5op2BkxA7aWxnWIC8Aob2wp1GE78C4OPnuI
uJkmfYeXanC40n0bqRUFgXc0YKvd+AbDZraI1T2z1g+732WbQP+7OjWvmN9tiQJoEF6XL1gjsV8M
5+QZUtw4FSqAZYL4kGf2yg/pAdSi0zaVhjqQ8G8tpkU0BJ55mXViatQ7FPO6DY3dXsFf5SIbWj2d
bZxuvy+WQIGM5ILiqtGBsj4ArgPO7k8TfwzdqU6nDVSUKfx/FFjEdTmtj24wdt4NMFw6R0gTFTcE
l9DMh1pITPmRuoDxB1ZAbjLu1y7Pw5lENpGgdrs4ETunWKNAWoWxUnpLAb4Nr+V/vQvIAbIIX9vn
kyy0bx6QejP6Z8zYwSgmdL3Nt0pMoShFHoH9Xc7xUYZUN6Q4yzgJm/ToXS7rNpKTGjbJyUe2Xpyc
UP6oPVFZHUK/nlkkZ7xZPCKoNwz1cv3vFyVA6GOjGrXb5F1Inf+Mf+FX/KLCKlRNJLAPS6IaLS1M
WUl4SFOH9YwjfDjnWCx7DnD0EncKWW+GXUe23YsagoSigu8q9KLCycN6tXjtZJnheSN/h5KIDjkZ
6W7Xuf8hR7IIJtGcSY2O7EhaKqoEMQrxtDERioJ2V18wOOmP6EGdcTLpVyNSyOy04Q69gSz0HF27
QDUL0ywsor8HB6IxnypCO6l9pxpiXFwR35RFhk+J5SCp/C62hQvBlp+C/l29lyncy9V26yMwTFrl
mlzaq2nCf3iWvURWBCZ+P6QFULRGbr4DVqcQDCPRGkfmWr4QcaB+fgL7NaQCnhSLx4PHHheuYuvW
NW2BmiqcB7SrmPsaKnMle6zC4DRBOJCj90/6gRgBTwEk6FznLLxHmyB4S6PI2iWc2qPP0d182kAS
g94/95KgKNzRfy/HA8jz/FtbFR8Ck2ElqiIYLJP5SpiSHC9lr52OtmJpEQS7UtiEFR1AFcK5W0yo
IeaDRXP65l3Y3VUQ6tH1PUloIKkwUolJAb6N9yXlu4CIEzuSXh0lbz6dCaHAu29pUl99/oNYHHuW
URjhMvbS4yNcj5jIzYfv6u2t1wppagCjzpN+FfG5x7ohxU+YTPBIn2K3rz76xGipkvxLbzj+xNg4
BklyqS8ghoTMxIr4NZAUOodUrPMzN451HsjuhLh9ViasyixE89vQq7x3c7DXuyGHRGsRbQcwzGnF
PxXQmHq4FvaF+xlsGwcA74lOgwdpf90aJIDmy4BrsFGcEYI28K1WXmxhFDiQk+zoVOp/OHHQXUvg
3aEG6aqpgt11NOyuepOFXnUGt4by2giIZTYQqe6uxIJX8wL5TNxPVyzkQ600adpQ/nwFW6LhQAu7
W5fHncjJThrr1hpptJaDTRPaGjeRn6OS/AKAJbdLfwFQ6bTUSrXdeuAarWRWLIO2TbRg/qAzWXYR
O0UMCGg5R52RTowcnKi11jKhVra8WjyNKs6Kohc3ozhoPCvkufD0zykcAVq1AXCIQB1FliqeZ/qV
0MvZMpCPN7+7400GJy5Q3tk3JcJxHiVWnq3PGIr8Rb6HZJQ1mwsO60jyrKaaK3c1vf2R8sBsprZf
ENRyksBBHXvj4Y5iCo4jI0ERGpjoQZBkdI7K2m7hEYYOU5TOVGrprtgxlYwAWoGuCQZZiKjkbVpp
zOls6mIvHW2elBdI30k8ilcQ23DgljgnZClL3/nFf0KLyGM/HMPtbSSdi238PZARjrdTqTNrTdVa
SE3ZmXH2Lr6DE89eRaOp/ZEhYnH0nX8+msm6lJS7NzzgzK1sJbW48bH9B2gn4XrfK36oDc+4pi8M
QqZvLR+zrqc4OodYGHTKqk7TcIDqC+PYG+IDNP1OoqbAkZUK2nRN0uhcIYEggqxVmRSyvfpYke5u
V267yntKXVrDgmpSRezTdQxmPCTRukyMPG75AYy/JJocsX40LNGpi2hpJg2GwOyEP2W8M5b+bRdA
7tP41/0MDD/U+C/6o4Oq7n69H60oZRNwyjrS/TNuJP28oy6RhbQLdcobFf4EZ2aVK5+RGhpKAtmT
5MmLz1bWJfabB3lIvr0EWkdF1EIVpv+MOG4q9YKlkox9xhzmB+pMohAsh5Dc2hEh0stTM1vCZjLC
G8YfdQ3ydxVjcurQCTBi3nRUlG2vznNMZKfSoh++doEuD/ZXv7FnOgX+pYOvU3yfzhL0POvI5vYW
ma8zH+0SMeDjq+PguG3giBZTTaD7NsKz3nMbmSDz2KZHlnx5y1tjl015tSISWleL0HlqnLmDr/MF
ItDG/MTNHqvMiEmnmvgpLnifl84/J581lFb+SxEvDX60FR4uv7iJe91VkPndxOJeQjwiWSlg0Jq6
Otep1it/mED157t08yEHMAqBYjemtaAxjdptKEi/dGoXh0HY1pADI3hoyMwN+5TO3ik/I4YnNYQ2
ONKgpKehe4uexCi8hop9S6bqGqP0Md3iDxPQv8//dZyJ0TaeBhiVQicnvVYehjVnBgqX+zIPRHZ1
KZZyldMqGjukmR+JUxBg52OUESQurQhB3H5T9y5VxqyxtVnIi2otUfmTLeBVDlHnbmol1CwyTo3A
AZ3/BV4LR03UyWDt/u0rIU5tpL8oEO72lFL0D/J0XxOMuDD90odIAumAONtR8XfxsU+uokGsqvkQ
AyqMQh/wkGiKS5KQf42rbG/Psz/wwPrwP/S4Zk5dZWZxt6SSD1jdaQXcEGIqULy/SYN6How/5Ru+
g8THzA5ZDLKQ+aa2SS7w8x4E0MRslF0EMsb0D1JEyha2ZQnAGBd79Ez/YvuvknMecfxefJyexI/M
kKCnr/szSSToY2sUnTEUyFKc8et5picC3zwzguLhJN7pdjrMX+zA5e6j03SKjTyQZYL1C8WY8RV3
ygVsFazDFx7MGtHcmQMPSzIh+pCwGtEO88ryaIu5v6sr+yK+o6rxMoGgpFtPwDcob7zMwutI+G24
4xEpRASp7ud96iChUsu6bSQb+y+PClMHMdseqRk0eVxnXl5RyDbzc3mwZlmY1OrSErE5I/NkiV7v
YN3qbe5C+0UsPZXreuMCLTptcyJkWen9fMeD81nNIxx8Wr88XjUUvCLDgZdlHA0VFYVfhpu2QSyx
2vP6qCRurDMnOFMFb1qy2dSt0pd7lDJyVJmrH74ePiKzCTlIE1lT/BDD7AaqeWhB/cdI8cD6ShLM
OynL7hc10TNoC0ruvimlAOuqlsGi9oRAFdZH25T4KMG3E8wScJ4tjRXwgsLIZlrrIJpGez+1T+Tn
hfwALewDJfM6FN80w28dJM3QlNMxmMsgtdJafXQU6foBct/Jl5CBksTSK0ZY7ryWmXRVnEVg3Ov6
ttvSdcG74qhp8H0bKBMKqvM8J/bGC+WSZNYn5AgnugUMSQfqseVUK7oHszOG2FyGgJFOpamtLFx9
MYloQplEMT3oKcSP6Kn+fF2NqVtvHnZ//cdEY2Ibfa5yeBmXy/xf4Ab2eagVYtDD3ty+utHPw52s
OLilvBEmmFvCryK7GRrckuMInQHvvTq5RQxPDL06nG7DmqcKt5Kr+AY1jW5AA1Ax5N0vUubrtkgu
tNomvTAZ462iDftjE/h7Nv/OxD8CuYow57VhzgWtlykqpbCKraYweRBDD2OTZgQJ72RlloCBhaBX
J/3NSPp95XTvWCJ5vwD4BbUei8k3bd2hsLy+XJmKNI3h5iV1UJoZUgsrV0Pf0eY9IHTwI9U/hqXM
yP88QBrL4T+y+ttgiUklfuzs3o5u4Mw65gLBAazbwXTpuGwCnFYxwHlUKUrKqjPRHFeM0Iqwd6wR
4zOYqgylYA5MAEJXVTExlzM/WSCUD8qLJskGfWNzck1ZzmFIgmtgNGhvFD2hBN8QiSLP16+t+0fr
tQpLc1wVkDxnw1ilOP1KRFshFJr97XZQjXdfQuKTQnrSpLrWwYZ5ZbhtxfazpqiM5AbP8lwnr3l0
9xjQOynhkPU0gUeO+c6GjxX2VO7L4cepIulgI3XJ2+hh2uNyVIVVHDghTy2UxNRpViVzL6KZdBWt
BV0yp1G/XAv1/EiFUuBEApd/1OMq6y0P2DCuj35+owssYG6B937aF7w7e/eE7M0lpvHCJsllFsFg
dhRuywbB0D65I53oferHeAo0l6wuyuJ42MbHMI1ICmb4yktdgvPPK1e2iGF9NAtxQmPMFblSEgbD
LOJ4zgTZBM7IB0h5IUM4itYuzjjfCm1HB7LrZo4rG1KUHaLazIlSK/Hs9Tgv/kro82dqSTR9Xe6h
7dvR8bYQUBBeIK5p1hyh0xt3BZxGYDdzutQDvhjhDxZQ+go/ZIssRrDPLuuc3au/AJXfdMljqssl
OEoofQohyy4x+HBWJkdK7VvSqKFJvwQcerGh/bPidAVP/M0u06qIfMX22mveiPCgFlZZsBJGXTfJ
NX5ltXClyVommSzdS5yOG7AcRIbmNuRGf1/O4jaG5OBBFPZ/sEyRc2+enYS4lmwcdNCl3l0y+pTW
GaprDCNZHH12lfTDRb2BW1NcIGRXRi2WhbcrYNHSpptJI6mWiVL30tPn0Pc66V7ZwCFafBTo8+F1
0szynb5VMC7y/xqgF99PlmKEV8AI6eVx4E9NAUwHTJDuEnnSgqxxM9EAl1ds+Z+sICwX30LdVfh4
UaSoZ8AcKLrJboRTWmlar+VyhnKrX53SQdn3OGrq64wyNgsV/EVwWwEHpOGaJhS1bwMd4ozlviVL
mv3lMzzFPcQg4uZ/RJ1bui0lPBMJdF5aPQKiLPfZlfotLcZTSsJflIajReyPyuYUy6qg4vAroi5z
/swda9Qh8i7Bxqf+nMoSOI6Fzl31V8Q3arg0kOUYfLN0E74VmdsmLPBNpQoneW8iR8MhJRm5lMSP
W2Q4DLGIfHO9MyhAbLtp9wLQ7br6ktINlXCIjiNBr+01T8OAR5R3vShjcgS1sOCYC9dNt9FF+40/
QkkWBIM72eQIvtS7D5xVF93+9fGu+zDEmbbYPJKnBS6sh7XbmfsgKpprRxW9iWgpD5Fc6a7Vk8zL
yRbvQptzIsiDgUtM0Bk1hZZvo8Zx43w0OyE7YasZz5TPLCr3TV/3CeNnF9RcOzbX3iaIrEzwZO+9
GQ2FDYDWCrXWWHzdvjTrd8nnxwI5ScqOCSVKWQhqiB+Sw18nOSxdEmLLoHJ1Cz9x+pCooCwxq7eY
F6SAhAkgWoC4TsNA2R89FAEmoFJy/Idkx2Uca+chdivundB2W5D124+OS7R01IKzAmTHOlFSapkD
jzLt08vP/R4lMfbcG5BPCy9JjW1PmuLuS6Di0VzWLlcFsVGC2d9uNuxwuTTqEOuJumf5eH6aaon+
RtBp8JF7JB76nrM54123N2W8/zw+GuT61ZyVT5hGx4MTgrZD+LnrAOmLkqn0dxjF9lvjYpe54prR
hRPLvLDkoy0TkYPcMcQwy5nLgpQ+QxutSVAkMC7wggxnzqZm8YlXHRsZiqpDPIEhIb2B9SX+AJGm
1oZ8gvdsExEs/h53vdKtXF6/WMb3cx93g+2jwTIJDVXqE0iADkIOBRSEu5S+NrTNLYxJvY128SBm
ScLeZ3dlLcBXT6pq/u5rVEupIr0TsfS0YK2y6SdrXWE3dVOYw3tCfmPvQuKY4Vf4vnXWtiJims01
+H8zpP/ZP/P2kYTaLcsrc+kIZPY88yTJqFdAur7ghouRBCCRJcpPxqxMPF7aH3grdFP0I5xpBHZ1
hQQT7Hp0pCHgU1u6IxDmLheDExWeRu4KIg8JAMVeOzFwkxZ+vzv7EIaPP8OPKPNGsjfzjlt5stWY
+UvW2JetUqKnNuF56zEtBMjqSNTEJUf1yZLrFNfdJDoZGaRCPBx1bjYQsONlU+Xfu5F3pOLRzwaz
mMo5D797daOQRii3g9lwAoppDe0CvbY/44yOJHTdI+okFO0jEc6Ge3eP6KffcYIxl525Pv+V9ZaX
AIHs3KK18ELTxJSCZOTeYWjHgAy7IK6W8dCLbqjxapA5BDIUJXgY5BnLDoMVd4U+CstP17ZNvmkc
Wis1BNlUJSZyM/aQnDgVjbtKSDYqkj0Pl8InbswGGnhIytTTPscUI+qgVro0kanuP68zNmE6HgQT
bQR4hyTDbwBuQQevgZdGq6P2bcp73m5UgLQbpSPkEm6MsHmkBam94yqr9YEEsIOtW690JGNBHiXb
UVgdeuX5aKcZncHyR5jxVUeiD4VrTZQyl79Ep/L4/eFTfCZCRfNFfbJSHjJZhxpmoSiUiNv4+sKw
OADE8beuCJbG/XpXRINHaKnDRVWk73/YMT6Eyt0KPlS5nTTivxNCAWW0/3BLY3f/jZ1DJg6POBn7
bZmDfQ8K3aMaB0qtlMSwAfJkJXBj0Oz1l263hIV9YjJ+q6XysImkWU+0yaGv7sPz0BNgeWPU8JRt
3PUQ7d0egI66Q1sIhufIFZJkYTdPxC26IA1JHQTa/B6A3mZ7X28oOCN+WBBuiSq8eRhk5ZRGALRv
6MrA8ax623CBcw/ja1GrjlgyQojlxoDBX2VThAxWkk10WWplEWWxwPTcQpbM07gBcxyG6speGfmc
fHnX9nXRoO7iZ36lwhglO2CbEuP+/yYZUwLMgLYvVsRYvJmEn7gwOa75ScGEzzOntM6VsV6/4ods
q5RU24l+kuuQUgDWKPMGueqOdvr76UOazq261R86FOoa5rp3aFci3rtyO0OgtsrejUkLfarwMFVG
ZxCbl/REr3A06/QjJEJL/mb0Dwq9Gjoc3VTz+R7I6QGc4OAia/QROU07cHxQmjAN7t+2kt+Bljyg
JUFteiJozkwmSs0IH+NsnXHPgwKOAbGKOLYzApEl6OhHVWiS28fuyP1diQMBQh73GwiEldc1q+zu
/baoC76Z3WPVySmdfH7Lp7RCe1fHziFYU/qG2TrEQm7PLrI+ccVY0jsHpZhzavI7C4w7o2+L3oFZ
nyMjybK8Ey+Iow5j77x3fIWiCQ4qteDZ2Yl6qPWsVBN695jRIAd1nQTKqoqCiuchrdlKwBtLl1AW
+G0vup5hQpHaFyjJQFBhmk1ExrXnuy0sBbZkPwQWqmWfbPwaPXhlwIFztQS7pIs3CYooGdmIeIca
sMTcfjUPUWQsrD7/qgsB8iqeFY/i8lC7KyhDf2NJ787huaeZ41XTWYs4jWvzpVrhWpnBpvouvfot
ZXWeTfjo6q3W5uMjecueGh5rf27vzM5kS4gAD906TraoppWOIGAR+4MjjyyqNN/X4my5VFAWPHDa
2lqLqnBvwuzRlukT+jRDlO+O2AZrW3HDCPaQXFAmpXrFbKz77mtk8FFhKlHJ6kEngLlWVHe5qLKy
Xhqpqf8Q4vdqQVbAhw68TYmw4EdE46yr/fgApoiLa+0MqhRv6X9VlvA64IpKw1A7cvOlUqbfo4CL
Hx3dQ28xaiU9FK4NEcGIhB8hPmAHHTjJaQDXEvXavlT389pSXF5PEMjfKt6EUcTbAIXvT4aPrIBD
sl2plyW09B2UmIkVr0C6ECYGCdaNEztWAk5SeU2b3nUByxRGBEMrS2p4qbkjh0Okh6y5EQ0ou/iL
FGOc4jPgV1mD3pGDL2cQeLsndliMRbcP6En60WmJW81LNW/XTF8+ujIFMCWg8QD2pB4XP2piIt8f
TyFkz2HPfYpbUiDu2RHlfQbLkiZ8N57a7emaG77wW4l3Qn2SUmEDASSNpeBZeuqBRdLErSSOSGtv
1d+iKQUBOELkD+OqBsPJkvGhgd1B416g0GX8ZOlSAmC3mMbUdHpJfW9SnjObe28qYuuIQB7us51Y
9ccs28Z+Y4//T8czSFga8VvrfWITqn5v5Hh6l0gniK6UjCtG2TJPx3En019WT+8bVkuTify4yLQh
/TVgJNFy1xTpCyBaazjNP+Uj7CxHUFcGMQ1Xp8qcoVeJsK6Trr1GBRhiFH4ogMbDewaoBDeUjoPv
oyzURqX8qoKChaB25KgEdqcimviwgHL1Gx6jjCtkkLaxvPRVYInmtl44bTiKbpLk7tRU8X5t2Tl/
dNd9OT3nQylDPinMNtdSmGErWwHwii7z0GQgioW90l/G4Ig+siElD0j+GzyO+rsBOhVysSGQUlUS
fql00jElDJCozNBDo9VM75vYyqURq1hMQWE0dta1MQVcobYbTrOeJ+EES0uLINz6HDMlpqYjl1eT
H3YQ6IVx/ngA5AiBsMjedsBsoaYyDnx+oq46Wcw4TRkoJJH6JdQjhUkha6GvxyUenViqyRQhFYGN
pggJrzPDPHe/ZiuBXV4hvCQYLNmwPnspiypuv8FNHTPDp6GN7J6Y7cEpsfzN46jcP1Q4NGUnaFeq
ZG2iLrlFTNfZOkKnIn++Gx2K4buGGQt4H7KD7ZwHE7nKD1SYKH5raUoXXce8dzDxNoNWgRBh5T9F
e6l4K1ko9nQ839sd2KiggcxTMo6+J4mdO6z06bWHuy+FE+NW0B1yKv1cicOb8J3krMi6CssIH3tx
7V0enAN3JlvQV0A9hPC77BO03WnhTfz+NFnD5aqDDjHzpDHLsPiVF4E4pW8nlxcP/pYxoR4q1DJ9
DxKJ41A8Hp4LnhRSPf97k3ODGi6BJcbFFnqCLwnh8bW0l5EpqgJGguXi16IikNcXvXxtgNidLzek
WHlL0hrNVGQkJjS/l84Pq7zG2i+En3ve1AsaKPYnlnLd5kS5uKf5KP2S7gXzco8049fSwMbKvmxP
4cx3zVpsVonuezoZ1XT+NVx6EwRHiZ434FAZ99v50NjxQMHIMzKd57NBMMG4SHQ/lETocxPX6orJ
4d0H9E42fnuaruLOw2OEV5S7vu9+yrCkFwz0BG4/WMpGVfgINTRd34CY0tfQHBn7rbi/q5aTxRrT
lF4R3hLyCbepz2ALMwxwRwjuZhM5rzkzdI03X5OIUvA9ElaEJEegXrBendIHgZwriU8a/f96hHKP
lx+MYE1dcfKP/zPa7DtjwEq321/x0KhP6eutQfqcSopq9WuOGomFcSl50lvluMXhEQE2obxM8YCH
rDivZFRZ+a02w73GZhpKyegccsKz4o4xRi+6yaw2AGbEZP07Rs+nqr575eUHPdb+mXhUZGkTnAWy
P7dgpfKnsneCGRPF5ziuIs2wOf6vEQbzSJR0StAHsI4h3kpDbtG5avr0LvBPIwL/U90c4/HvTy4Y
hckYi9qP+5BJ9lTZOEJnXrbTzMclR8ImIZN0TG8lVRc/7HvZ/hRtX8tofhjUjyMlJrt0GnAsMTLX
6/CrbTVB7jbbbDFkWy5WoYzLMt/YOmCAVcaj0iUDkfXdb92oeDwaTp2dIcNt21NGJgBXkl4dcdt8
pvT9jbybtd4n/s7raPIHti5sAe8pWVHDN75TTyl0rY+BK0lf5si7UFZr+eIlHqNq9mgDKPj1cIEh
9LLKVzmnXxePB4Es2uBNXM+TLzTZyPnqqF8R3JKr56Kj9jQDSmQobJPirnvObMAzA8tae8BH7jg0
VA3gjqwoBb3CsKfjPmy4fQWr3QiUzv3Y1Ru7/Gorw9FoUhURMXZpY31jnwCVD/LLeQQuw7jICF14
BKY9aG9CZFZqUYtVfupKfFD6jnPCiAcbov5AyymTEO5RLRoMcW9472/ecKTwF+FgLO15TeLdRWSK
uftUNAtJC7sDFG0H/1fV5xB92zyVvjrCxUiYmL/rAe9MWbcSc39ov0d8BAId4E2XXK43ir3dlDC3
booFAybDy/p1R2nf/keSRmmuR88fqNAmNwuxOnvBg2i+X7pUFw7rCtRzDA6S6fbjsOBn5/EIe2sK
9lbbe10w3XHjkEpkIrWClFvjN6y3kE8PRJejtz5DhGqct80BChOAG4bpvSBfD/UhocZd6TL1zAEs
NOe5ApouCimEVe1a7Ix/P0wtu3ltmogDhta3jbia+sX1KwsxVQBUSxhhryMkY8dHFJA2BuhAF60v
4Hi6eET7qaqAFz8vcQNPRg/1JLd97wnOByf69Tx9YSYemPCAF1fQYD+l2Rj4fapChknfGw/uvi/S
r8+yXNRI4xmCE1FA/+JK71EcivEv54TLbM+Uo38gA/jvfgNxa3MKyIsqHlIwZ92o68lWG/7rGlqK
XMg7jFBqrESr3jHNfD4v1eOwR9TJ5NNNvTRQNVuqU/SBhtaQzMlHZf8DlnclUqQKiqQmsNdGFiDP
VZiP90n6eo06Ut3IrGYzmU6HOZRAsSjscVHfzBTrPi75hVPIIPno4boOB5O28vBIACvguy8lgGBA
B/Cma+KRbbvQrNnnoTcTBiNYRneDJrAwJEM28tOMum4zLTjqn9SOJjhwpP1M+4W8qFbHUCC1oCgN
SX0ImTLA6NUWK0BuPzNNsa7aMqKnUBwGlAkmOmZctEuTNksq4kqd0H1nuDtpciNSuT4g84gZXg5s
glZEIWorSAbHJyoYZdLweX2Zc3uR3MiXUzKKJpMcET4W57MKvgu7cpXKqAkrM40Wli7D1mthuGYy
ZPWvBZtKWpfNQD6f3dL6XYbnHfegVYubTb2ZN59+Q5jOrKMEg36NC3ewF5x/GlXmHtSeuAfB37Ii
8ARV7J4daL1Z21KkZdP1ncr8paLcTV/XOx/IPXZIwddnus1y7Lc+JK+PSqzvW0mk3iZD95J5eQc8
WFxXVxjDNWvozFNIrUsT96XVo/BZD5MNIhyD9moXumC5OLktd8el6lB+djmfIrdFl8Sli2QGVhdq
BVTEvqG/WHDAK/MwcKaPmS8UUYIEqECsb1re8Yi/aeRIsXccK7ZdMogOz7EPR0J7/liBGSw1Jf54
DrIuGEdQ8w6jbSZYGhTQZ0QUs3s9sC3TpB20er2P+po33b9HZa+SrIJ3T/12GwWTnWRl6UUlV9IA
NOpl9c2VEwnulF0LfTQMgwhvDhVx7+W4fl3ViYggJCj8341vXbLkrOLDmTfSkVA+XKHLMRR+euNh
poraIrSJgQHJkpizSObPyJSnDGzgyjPib8s1Wl82FYhFOR3Eu2Ic6lQR4t4owtrGwTBwcVCuOstg
hA6ula8NlhnFoOLj60QqmaS79Yk73hUVdFOPhDZ6e8wdvfa+xHr7tvw7x5ol48T3wAf0pPPvEDhh
YTZ0pI9Uv3N0KKKjCEDQtfyVK/zKvbWARcTu8HQZ/EIRCEfMKNMGnwOibuYHv3hOwBcyPhbUZx/e
ouHF0vHcs0k3QiCLpNzXv5g7xaEck/2p3ZiiRwY4w+nxS9l705SplcAN+wQZwnQTW7WywUax0Hif
U+t3C9Cm6rgTZJv/P++CiCN9JEzE3+Zke66LmFRSC13AlHOezxJGqpzbz8czwA9xeWVstsfvdFy7
fOj2mnu6gZW8UIkCZ4lcrVw4K6WYT10i1418dnLnI0qQ7QNy9fKYgn1dc37xodUsSpTZg7DSHXB2
uls0Fas0tVg+TvpNPUiex1gwnggVJXvzokDGmazgBcytsvQlgJB58YadJmWHSEhhzop8COolecde
2yAaWzbV1FhWKkSlZboppXlYM12rRCVTVMxir1OSIJT9dGUyYg5T06Tm15iYxAYDShZOPehO1ja4
QYmf1A81vaK6Rw0/n05jLWH/RQE3An87/LSAo7g6De6AiVGnu0IEpODGNg4tl0iroToxTUSRHP7G
Zd8ax7DtRwqFmmw1zrXU6NEl6sjsh+O1vP1+ZUKWHtbtyFBlWAKgQlxDS5E09tcVQsxmcjKxlTXa
8Qj3cCELeWrizkYil1j8L3Tla854fm7wt8FQ1CDkE9ZBqUSl9iriaRI/AgCcgzslT40ToYuwqZXc
dez0XCQCYjTLjH1ugUJIn6dmy9qItxDYrHIhuwU33qVwf97kGtwGZnXsp0XwKnwR2sH+oqdpkgAi
/7Xk3yUqQ8648SjXBIF+qvbl9iZDtR5pOnxDaNNnxCOr4nC5Cm20IyNdLkmWhtwIQIXxPbK6y53x
iCIbvcKjZbZhbnG4S+vAXoR0iUWm309FakdqUOhN850mBfb1pg5ib9nZXXAm7LLgFzm76T1BdDCb
LguAnPLhhJlaYNJTsBduZj58orwPO8JTa6oQolZerri/yRpB5gt/YF1KHdTwpL78aAtsrvvNseC+
AWpf17qDrBZpvMIooX5sEMqdshNgIGWU7dtgZTwxSuxa1v+ZYl3xkfLm8u8yb+8cpzGUK/SSD2bU
alzNRz7jCXziY5agYz90ioPmcUBwjDDgdaWPhFy8egYQbLREPnqJ34C+78ikLVFxw87OkhbJlGIC
eZ1g3hNGH+eSJwNFKRNrC9tbp5sZ4Z6TX4FKXTAOLy82tTsfEJW6odAUSSMzxdstlcekOQTe/g4y
KSuCNzhQN8MA5OhxoSZFzmX9F5W/PzASnpMF1G3VVMbN6viMOxixImqBWcsq2PI46J5M1BLkt2XL
Ny6GXeZKKTFDnXuFX+m+vtmBbGngjjdzmFOhQ3CPFxqEygmUTd/9oUyPqEcURQ/oa6N/wxvBccu0
nu8mYNeDwjyzkupPkr/RaKwymyfVwHVO5XNz5qhlT0c+GSoVLusr1jYXctITFxaq50VKobi5NT+b
WuAJZ8TZPqgEu+SLIg9Ar3NcM5Z0sWzqLuz3ZS/zC5PbReZYDkMGfdcS8O8GdZuQzGOUBmeJhqye
zI4DyfvwNY8LH6XeJGVkEnznvSJmcvlqKIqXytfxvX9Qc8aSgvY5we8/nN8qq975E+ecu9JhgeE9
wSwm2mQ7k+XW7/VhSZ3HpM4ZvkPmrcDnEEtN7PU05NjkqSU+oynb1Eu2ooQJKRBnyNy/D44d6qwv
FizMWV0rbUKh3rOUnYFsk2MMTOavViM5RhwhtVYYIQQh4WQsbW24zj/2NGXS/DynemkBn8z604yT
r2Ey9VgYNsYP03XHTztXXkJBPrrSApf2VpLuD/NnCvI/EY5K5SURr2B0+0eR4Su7bd2j9VYaLYYx
xNi/3ewuipvCD5NIa6v9XuvaHR7itxbh6F57fgtWQ0yrkNJySO3+6Q+11dtds92fMozIO2aFkU+3
GAUrcn+r5blNbnRJrJUejffctE7orcYG33iC2nRCk31vV8fyqtKf23c4WrgofbrqT7xL4Fv9opAf
0/zj5mZTOFFPSMum/64bu34QreNTQJ9JJd2wdp464eZj8etGYfzgmO2/hNAHllEQPVIGCW0JP4dk
mh2JhRnmYUrf/yJlvfp4E7Bq8KAqvAo7H0npZrLtFne8K1SqgYE4tyg5DiVxUWsCJs5wOT3PDV3X
2jOLQwe8UVJrmplL90YHDXwpcx+sOszyLVM6hQ0BQpjl/TzKKiYv1ug+shRyKpBEE/bam7KaI2hJ
1AoXaAYzOpa8/agFKAFgqLZoTb0yEaxDRr1y0u5FNi6WqKIGSqsywHuJChgxjWm48Y6wsxZxGtjQ
LbtdydfVOBwfdpBU6slmnQKKigSBU3nKAk8ii0qRQ3rux7582nJ1MHwc1AShvJjJlh6JajhWWuLI
cO6MHW1xS/twV7FVVatOpW4JQzuR6143vkmDT0Avg5rLBmniGAHnqzjVdqd9OD0MFy1Y9/Ye+U+T
JyMRrg8bvnb7KO3ZVvn6Re8lYFYo3XkkbcDOocHH7eRWZR0vaV+lij5nzx0ya3HcULMLVLT76yAS
ZtKmqpPS2o8nYTLQbKHmyUtXSmdDPVS+A+YK+tCDCpHrZG4P2EeqpdDnGeDCb4Vvy9cs3SC+eWAH
cSkrTMSnKmTWm434gr3AVbmAuuxfuYO6AT6oOmnzPJaSHJlDGgXzyFv2foNqsTDCIP3n0p3DKSGu
erqQGmH93YibAhH2Oph7x74hO+iQ+ZR2EhhlFCl27OQ3430JscQvWjRUGI63QS55wNFYrZWhZN2I
ymQq6QiMWpJyxPwGHVoc5ZAElp0umDPk7EviE7SqxgfVBZ0coBuXq0zbEjxAcF29stjaWwkjtdIg
kQnHzuedqOjObDnYJOjqI59dmSPD+a6JeoIQS8k5QIs2vWI4j9aQiJjGGnK8p8KCede516khhhi8
2BO4VWYAHtOdEWQ/x9oKvvFa/8Il8KaOop7yii5bnbUzICUXkYUgyMWTjnqFmZNeiqpXoaTrIf57
kFZNSEJMZav7QuOmzfHuZ6o6mUaCqcn/xloFfzmfQsdBK0NeZ2V6gC8WqwwXxWfZ+Dr4vWy95A0Z
eAAMGNIXUU92mAoXpUqw//M5gPxzm0FRwpC1/qfK4gQrdtIL0qiIfRmugk/VyJywySVarOzvLa9J
IB0/fvPIA7a5baCt8G2aO1ew1BuI1YsWo5T6gmgZzvLEfbLyOox8ZhEVmkxvmeCNjTMMqGxitbKg
Adm6teMJDkcYne7yMWbf3VI62PP4HRsWCto+k47Zw0zenBFqTbfXq6E8Rh+foLwBm5NdOkQJP9cR
mp2UKBqV65PNd82PqOBBqLh7V+OJZA7NFdzpgIq9TmVfJiPdeImSDLDfHxTHFq2TxF7fGs85sXJF
s3oRyQmbgRTeKv+ylf29EPgbi4Iwr9D20XnnVBz/Hk2Z94CpuT3GKiEThqh/vMGgBqZpqzbsP3R3
8iBG0qbJMisQJmtcVDvoa8X52Y1rhhXl8wLWaUeDhUX0yv7/yNOBD/4R2Hwo/G5qGX7Cxelg1hS7
Hn39UZzqvAqO0S0fuAnkz9clo6oB+eeLPlay/rxDU6EXy58trzcHE5ZC4MEjKag0uCdXfkC8GLKI
v5+TVOcK7Rq0di6sfXaVLPW8Vi+78YPD1Qxn/ImssoIUlUfH4G6tlgrDs3WAcQID+7/glgVUUezR
N5XH6ZmTIDICkysEvjY6QvMuzyIJtiHs0/J/HWpZfYJfYew1sAhbbEvl9P8y8WBqD+SNNlAaw4KF
mtZ0Gc6aMZ8OSpiil/ldGKPVvmCaaXa/D6fyYvGSiPCcqHpCV+2cj8AgeFuCl63SbT7d8vElQG6C
sp83KvRm17gYbBiM6anW6cdWK3oJiEGwHLpPMpNCBDxCBCIAUhuX5i9Db8codZXgMMBxoYCAk6h9
ScGrsQXeq4Kpw+od6lKyNkn0nl3p6swEfmZy8wjE2JoUm7IpFiu/qaM6HXF13rlCXlWrd9j7pmnr
N1VhuzCwwLkBoGX00qbuvhjxRVA2BFl+lQpwfVhfm+aY27EFt8u3SdKLV7ekGXy3E1akKMseT8oJ
Us1KlUsg+jTO4rPLlDE1h26znTr86A6YPqKxJHk4fM16nM9eAOAIiYGlZ5Lvbw/dNusZ6fYGcM4N
Vivqm1djaccsGD6uqAUZkRIxCzZDSc9lOIz5vyJD1kHd69L9Bv4oymxakFIA70ww5mscLK253OgR
d749cOTCPeGroU9l8VwiRgGwr0E3Wtxq+LzpTJ6FkNp3j27AA7xgv9Sraegl0FBOWIbO04+CaLtr
E40VEeM0pvowffgE6PUAW61NLCk31zC7k4OEiznatTjFfbAP/gpAMFDnqnu5Kd/Img31JiG1jImT
ja1jR7/qecnIg6uimyCxNudNGpnDXYEDTynigKuAcbdDuhLdtPth728+yjnXkR+c2RUhmsvMDahz
PERKneN2K66vXMI0wHdHPeUICWdket8c0PgfUwotUopphw7BkBybzhmEeGiF0snTBdu66LQEOXUX
Kqq9Ncvkvd72HuVtDKgF6BtiFj3wdf7UYahY9r9f9cPnQi1V6eGBodlI1IdFkkTiKK5g3ALnjdJl
VCSgF3Od+5n2b+FwjywgR8QzipYQPq6ENlqwcvl8Qjh4qugFgkw+qP0xJNI101J4SUIeIJltjmha
Y/bbCAlLVx24yZmLvcrD/DUhovlvew+W/H4MVoiRmA6Jqw1tea0jgohpM/3vbt1lOq62gozaPB/M
Rp2n+8/svR9UZtYU4LFcFMJUie1HCcztsKIC+RHCX/GG8gfcijizUacdpPFXTZ2Ybo/zJeEsjX22
xGJvdN6DKVuuWP9Qlf0gKZTrACA9H6YSclqmD99Ns9NXnxJ1xrAoD2l3QdbuiXQKeYZMXKsQybx/
CIYSk2JhWBF8ayQtih6AuJIOJl6eYRzBIaGSKwuyY5/r14GSih8p4sePGukBqWebQCxhICMJUQaQ
6vmjc325hoJ+2rZPVZD2OMzOIysUCtAMJutHjtlHRS+1gJTOV0ff/NTpIEm9C6oyszaZ0/VTDsz1
cPkjSi7YsEplZ70fHVh+eoJ5K1pbv9N0uSDz1SgGL44Mzn+pec5Z7zzJ9/NSjA0t7exx0KJVcfqI
0ekUIOLK4YViHj2H0FUnKPuxAewLHvNJEbLzMIa2Lm08Vkd6+Yiu57ovsu0KW7gsA0avftX3x4cn
FENeEndH7kV9QJY2J0aucTNnpIrWyniHaRATZnrMtJ1eVMJhFD+fTA7RADNbAO/E0Mvci2Va1af8
LFtd/5slSuUOVT4EljCb+kUSEUwiM13gOqgx9YknPtVSihRcppzqpZ+QZ+5dzLZ3UmGCaj3f/sUG
vMcrYXOnKYJRXuejuH+qK9i5LGKnclLwhROwbSAaA8bm6P3UyYN9zyoQk1DME6O5GvjJNWHKVA5x
QeesIxY6Xya4kTacqJaiXwk+WO0/aq1ByZoZkxNePdNVNPUe2wotFYvrUCMcn7zZuKUB9PVEVVyH
JcvehulHGCmWIGedC+Jna+4PMJS15JxRFQn+BL9+jI26H3jz0VgDeGg3b1e60/Cz0fsiMn4J6zrn
RsIvPyxwSYbAV+hGzrv5klthOQXiiQbB6h8BA3udhbbpd+UMQNJVRtyneoDoeb5Z/0WL94SxpYG+
PeHrweBrq1aN96n53XgfxI0+qkYhtiMNxSO7sX9k0Yb/cZe4O7iW/mFGYPY29K5BGgkazhac/LYq
5sR0GFnh8UgqJZqpALmsfA5SNyVJncKDNTIfORIOLiLnn85BkLDe5m03TpwaCfMQciVxT5jSkAHM
TeIdERokD8gFKVkGZyx8hky0HqEolamNVsNwyFtQ8QAzg2YBWORUhs24hr4zEIgKj/Esk3H6aJ3H
+M9u5X5UtdVV4MjzLpkPb+VW9+nX6hJhLMnnuAxuozKO/+yeTs6Gb/Bp0BFs1R8gU154BXsw8QEh
Nhnp3Cpp++STbq3NqSHh7N9j3RanKYFUizfpWE5KeFJKD3ov5zEHj+Vg7CB2YxP3XqLHCttNdCtK
q1pXSp9+t08ESEj5bbsEJDNlRStxOkAuMsxdwszyL3oskYnkJSH8oEG7mJ5dZWdzN675+7TH/yNP
OWPEwv/MQFkAVxVdbMflF2yofj+YkLyMep8aCY3ok66tpzFs4MsvBTrIK3RNyKGw4FswWQlWV30V
YdS5xpjhu8A13wsD1dQ2FX8p5PdpBJ6s+32N+Lin9ywJcYJmYqVd4Ieq18wC9dJMRpNjp3+dZnTg
zOB8ZejjCpCKo/c1ScwWtj+6JefL3vQQohJcYI2SkLmHrtSQ/0VQRkXlBzrW/2g5HadieHa8Ru8I
EhkTgdjjS9FW6nx7HUcC1qt8232L/d+TMlYkKD6XA5IdGTqENvq2/lZkZENwA+Y7+/7mbu28Kvkm
QRaTDt7rfDx6HEUI6cQWke2+llVDmOpyyMtMVqztiNqH30kwTUti2Bvrp7cNWUlzmg3zJny45NGR
2YlrWsKVVoh9w5eo8cZmelraQSk/jEmf5/Z5wkTwYtURz6J36SlNjFlX/QOrr/JjdC0S48A7Vy2n
XLlWs1ubB6zCClBwEz1KNUs1J9B2lUwhiZIrayc17ALLiEnCBW+iV06PH2NaQ6JPmlLDXVAHZkPw
h7Y6L5WKBMAP9ATKQBvhLCu7e0RxKHpYYtXmUBf+rPIZxet06Jm3T7HOmCG3KoJx9euBmlebwOD+
7zJyZj+93K8IZrwdU9zogPY+UxorYkJtGAoPVnhYEJGwgtYQuXZAl4j4r1W0dAJ5tLTTo9pTKKe7
Hen4WYQkmhoCuq4gNAXrqOlnC8iYYqRXka0Miq4pxIh+8FQrVqkEFsPPFz3wLPnX4ft3SLeamFuo
sf7EiPFh3lPEeqLRnMiRxjXpqADyl03HXRdpEx2rbpovyIixamPSzRe6CJXwzt58pYsh9H12s8Nf
iB4ZAM7WeLZo0bRouJL0puX7nfc3IdsPZ1r6bJYeo7WbETNncA8OkGBE2RIaFVScBifdVKz8lUZK
oeO1d25K3xwR+ioOEKxGOw//PT3YEDSfRLv3Gtw4Vo2lKbCI+k5oTHwnbEkhHB1GXmSWOMft5TqV
4RExllB1RGuxEPTWu7KG+yB5upN2PMDExJIQ5/kbzy9gYqsNwWwrLkL6rzIMqp88gY0ln3r85Abx
WDyrWDyvO0pim1U9NLh7AjtB0xYON2re/OgflBwlxcHwbL9s5XjefWxqi9oPj59H4IbbCuVhEuOr
9VOjzYA05zZBJmnWwCYeksVuPo7HQ2J6p9qkeUF9lUEaQVv2pRLfwR97dQvtW6sQngcRewdAl9l7
+KPgjQN+cjrEfF1i3lW+VWHDmy2J6nlFAxgYqPAWJvSzEfUfsFKXBIXciRLVebTBam0T53JI2Jxg
iKFpZWvnNeMWBM7oQ1K3Tcuh6iJa061QDDDI9UwJej7nFy7dgfR7XZPhj//OI+nSmoFW6JhrLJ0I
8YGXVPsVbbr0gnZzzFiYbxtO1r6/CQu+DLdsoOOszSI1MvcPuF51c9xTB0L5kn4E6dIyB3iiP2xh
zMLAH39b2EfVgKb6SbVOKcGU40Co7u141RYT4cTmPyunyuLiCwb/4tFm1fhDFxIwZDty1bOhyeW3
19fFnjdGt/DSMkgK4UjnuClyChSF/D1nt5UnGP6j4QMUcK5G7EfIiZL5JI090pYtDe2SGK9byPEv
SfoJyHUlp+DWwpdrlRo3HGVPHnbAz66uV5bBQZ4zQQ8Q5wIswb6XbjBoNsho+uz7w4X1SyE1nrAi
VnXRAwxgl4cU1YEhXQcKAhQm5QG1aDBEf+op/aZyz/IEojZSz6w1CSZcnbMmCoxpruzVLVd1OSFs
Sn8WsaHBWboxNOKBWbElD/bO/ShF0pXQLbopNaDmcQboEHdipml8qTs5B/gi9ewhxZB5JJmuIBvz
4ZlSaRCyrdZTkfdAdsekEUFg3DIj0Lf/adRWYhElCzUvOlXPjZmia4xr9bwER42HrDrQ3TQyrHDs
D6IkACtqU2cJUpe0EMJlVhJhlTWWc8AbBrROSpfTps+QA1Jw12Qc4HIOJ29ybgbvKOqK05dCklaS
rWKjNIa9oVEvcf5gTvoKZ2ozFl79TzAIrcqcabxVwbAXdNb8LGJpdbDTQPd8kbFJcj0hT00+dvBa
0Kf4QBBX+P4BWWdD6SwKEZyCbjvf95PV0Cs8r/gD2N3IHVwB0V856z8Irz3SFzqoQNqLAlmiyNmQ
sCBbCi4gsqrT9IWPuPD/C1VhwzMgxHUyY1sRiThwf+Hdz6dmIGNYkCrxU4Nd5Z4VtAn0sRHyiixU
ShSzSG2Y9bBflS4Jm/i96TrYUDYodCzzlOv5LRbqWzyHpmWVT8z1pgGRFT3QjmrzBS3ivfR7Oalz
74HpS7hT1ou66VVq1JRqAMepoTj+/XQXBbCfvWhQkrIQiPCAJFlXdn7Eh1nLpBYgJBd6rtp37h+D
fLzzMPqLCjcdmG8fv/IqNbGC4qC0zLC62vBwi0ALbetv0wyxUtP5XAWgyL4Y1eH+xZ52pBfiCE4v
PnPEJ2gFgteVgE21vgxFPNc+cs1GFNCLbHCRXIU5da6OOi9YJS31x8IdlOF+0+45RTmL3QDYy4U5
V6r7i8I/F62Za16Mml0+JT0Avfup+XFqgMR2Fb8+G+yPu0GD8kVAgEgM0RzBKBaynkJxIGy0cSdq
tqnxUBe8NBUBSkKXQmBa/+wslu51YPxLrkVjOLtlocRzJrBiTaWnA83CHRsfLiYaSMBLG+/42yGm
Z80XJ6ROPDcJHnXfhFHxws+BjUGTrX8BJ39AiR1/tyzz1dNXFTvqIIHEhCqa2w+ZLFNBIagphfls
cwt2CcX01VLYraJFLC7kfVF74qwaVaFaDjTSPzlziOZZr3cUsy/glJKX8kpOtRjsbQY8DPSY9Y7V
lys2pFoQZcf6hIY/HZeMndQvV0CHsIbENWQ0UKbgNY92xlMRaG8P9u8ujrq9gEo81s1zUlnfOuhm
JIjqiLq/sMExXmqfxzq+39hpgMjLi170huOZJiLOJ3azaBRICStLc5WWId1t1Is7NjNi8RhzNMPm
wkHdbEz47dj9VEpRS23Wd37yZp6b5ukqTuGq8nEWCg3Q5ATn+1O2W/Xq/AEdeZm/x+dNIpLavZb4
rRDqJjhadqqPEY7oRND6RWFVCHduira8g1oVNyR3MGjDFzZC7iKsAwbmKN44m9OHnQA0gXOdIt1j
kwtVrXjLDNdXH3upiqYmcSgTJ9vE08m8TMftjfQi5PJHj17OuXR6otVK8bBWvNL1v+pMieATkQHp
UYZGxSJy9XLBz6PT/v2Or5Wkbidr3BERaRLG7pQ9ZOvNMtEIQH/K9H9EwwnLOMQn426tgj5m0iRH
qTKs+d9TD8lYLckcivxixBt4OTUGY2aLhmnMA8eT691Ye0lwAJMRgJ9T/dLQ0VpE4++fSRWGheEQ
Hm6NpP5VVnwdOAQtB3TvvFZuK7HWJnnkM60OcZeX86Wu79WT/yVSHRCogUv4cXNbdjPJUnUkhDnd
trzJcLQmzbXMhV568isrkxLPU3AIItRp2DpFxXxqaMyE5vL91hgqCLmziFxiwF/mgffWoqcOu6wr
RggMdZCNmfjMzVP2WEDYRxs6no1kczSGoPotl0zmYAiMBlKc3FiR73TzBzCIv3584I+jVkwkCFqo
P6w9qHfD+qvOupDV5oWTz9lonqQvk458BGCbRaEHNgfBGUEDT5nfq3Wya73NQ99qr2aOqI9T5Bv5
Z5Y6v+LBanwIDQq4Qt58cTKbFa16vKzXuhvdoBOFuI6aH3tKF4ABedOleCkgLf5IqUicXtu/t4RL
FRsoY4hHAOM+2XreqLPzxnSNx/RJgtIh/M0P2KuJJG659TUcUN+MlGYyD8eUNwHlVWNOpHQ6LmSh
wdcRjYO/tJBgWhK5fAZbh+yKIm5E99z4HqfTjvihVmLftLclItpO5TC9XiD9JGiwHcK5QJT+RSpe
f8S/pobnI2L3ZXn8UAwFgBtRU57p+t4kczlUkCKIf1yiesWtoPke99bc7ShNqK+zgGTSGzpgw+QC
d9hveDxAppd9Gnjm2fbRZZs9DXq0KAXkufqWoqzzELTZufh6SmisJDOKB/DkHcQq6QkEMZ3rL00z
X/K7HALgaumA2No/Pkqn2jyrGbnJxAwWJQSvWsj0FQLu3CnvazafwtSbc9P3MR6hVzk6SFpypnXq
C3WXQE4aBKiGoIfIHg2WJ4ZBL9n+pn3aNwxmvjQgHtPwncvfTwlUM2RXjWeiykhnta+JBO5JsJG5
LIdHLAj+X+qvb4RSu9vDy5sLBCC0deY4F4aOiDoeUyQOYJR45LJfPshNj+O3hB485oUPeAXt/7l7
qdWYN8T/1+w2gl47Y9vJggtRWV+HM4hItuUiV7NEFPGY06wcSSWWNRdPUNbB9tCnxqujRBBCj0BE
CydXIo3clMkFjyo7AFNU+erBiXFTllUgJFB4MYawv6NW4Dsqv91DDiRs6H/iic6ph8RQVMHW3dLj
x+01nFxjDwvtG0MeQUXYDlwZnxpsMMrRoOelb155gvQ9TzxLxj4EfdtyoRWZiU/ExI5XXoBS0g6t
Lm7ME6Qv3377aS2qci3T0OKRHHJXD9PVGg3XrsOH54NRHQq5AzUdZ7Wbzh5vQmtHhb6mzsU4fFzD
h0+oWVcWrrdnlHGxUdLd/SYRIGqWWdVExxEmL3yu2TaTEcGZvAKgGkxDPvo3OiDtB1B0Fa76UuSU
iqoOiz35K7CSRbxQkDYbdwgjZ/LlgTdJpTo1OUXgI1qJRF70SzoCKmvWWrunQTJD80SBT1ffL5hL
rR1knHMJJwUm/knVXsOh67+dHb8GOb5R+SkOOOLULyGdoj1Vt8KLLS+q4ouDz+Lv5hAX7UuEkz9s
FGC7Y1EWYtZ/Lctja1c4AiiVFonfprnXe9Lqud3EHnGkiy5kTLeqduDFnPQbOzSoXiPOHIDXkO3E
cunuaxxLq0N7q6oezbof1uuDSqZADhX7BGndOmxUe/ij66VCIYVCMgvj3QGxIyznlvYgJewJ0cEY
C0WuPZjqhr1gv1yQmMCxX6XE2ZkGGCf5uNtMNZNxOFsE9Fobj9NtuAjfp8fczvdzkcm0//fSRfhi
1NSP4nQi4d23T3FSLbwMSeyWnisMjCjKiTf8urHouP/VZ1JZ0hQJ/xmieHA+iHDD3ZZAYYdGe2Ch
Bpuf14FzdPZvlD6Zpju/IU1L0wUx4L/6Hpzghr/PKGvZgE8U38dyVS07QFtm7zfHsQAXD3+bJm2b
Ewer48BKTQe7GSOZQ4mAFqpZCqBNkSZVCRe0csgOct76DQSVMd2HKMiAu3cN3+66Ynx/ZB9Xg7PR
GQ96so824vLdYcA+aKTYraLa8mP08bkGc8c/xHQb7v0/SKpD072G5W76ftOHzUak73rNgFx7oITl
QPp0jDEg7kthOwvaIHEKf/IG0V1GeLgO6p8QBqeIbdZd2ix/Z3Gt8LpeBT6DeI0iceblj30h04KP
lCdx1wGzpnk/dg85kcSECxGewTaEJATMo2tIrrfR+uB2ypGRsq8c9lVpVha0msXAHpIpO5vuxxh7
KjZ3FwFODiakho6wQ9LC+6vbOB4xYglw/G8lCDKB482FEvx2rD9C78d+qvQGopfTxddkvFxZW3LL
w5AVM2novnLi+f40wZrahq5ykZl+PE1/0d8mJwzQqYEZSHqB88e2/Rr95xpO0DMhOKZId/n4KuHh
Qf9T2SdH9n0QuyurdrhEanH9JU1/14FsknPOzayLYDIcDZgZWY8IUBoJqc8/kUE6kKKeIb2eo1XL
ccr8s/M51jB24qPHlawfeY35acqbIQ9XbcVyBW8XqWrnGN9QibeG0v/Z528TpyeO39UhR5P7FQt8
x7bnPzCIV2yOkfmkZMDogLVP1w/CEWQmNNTpDAbzTWsxHrMLPKBRWqE5u18ufMQBuLtNlAMXJaNU
d/TuNdskRK4b2/MTb5SsgYZzPbz59nqdQZfV0g7o5T5vanH669XebC5pbhL7igGyJxinwILL1YMm
tAxfq2hfxUhXyIdjKRLmSoGV4GEWN6+p+yhMKKD7zBvaSGN9AFWoSGVgC5g9jWFA9tNcOYbXWc4i
nKVU/5rx9hfsFwre3byHgAwC8DogH5V25se4fZ8+/YezA6kyEBUTKTQGGUcShYb+NJMBOj8N7UpO
iNSnGDGRAicr1ym88cbksLWxq+4h+fUHul6kJpR4iwkKSGGXd/OSclQQ7aWfladR777SrhQZUKL/
R0KVrSCmTRJ0dKqxRJ4eM0agoUMsxxyEmte3KPoAAU9+XR0biUy3jEofMKZGnbAiaRYbSE3RtbAc
WUBUX/lYQbc6qOiutEaXS3AA6whZmedsfjQd0iJutrrO3q6zi0qCcK10L3ermR6rhOfGKhLUHwvo
Z5/7FKlvDz+KpOeGkaoIY68PlHuQgsUmcfVyXVKo9Na7KK5pPuM1ij+EeHnF6KevI2KCEK1jVPUV
WkBcIzII3DhbXWFctfVXnnSD/CsYNJcV7B+PMXT2QDWYihbKKjS/2vslCg3XLTd8Dh4VjDtaIxzf
A4Pr1Qz03pkjNqNl3/23/hl8uT9lxDNoaFk3sILIAbcHpIX6D59v7MsMhlaYBnSqXNc5F5ivR05Y
7Pq86kMA+zwCEJzBMTGBAypeCZxnHkKaRfV8aKWSosJgrWjTo+u14WmAZ2T+zsgIGNDld+cpmTWw
nYcz+civd9hIvngGzOYFVzIVIJOjb9hpAOZaLWzya53FO7nQ5RS+8lRxtEeBo6us56hLledbqkWF
NnVtl/O3Nqc2fgnlMB07uG72DESElQlSC+4KQJTW4vx3rUTBBQs4fmqBrDFMwJPZ2XcrS50LSA/D
qZ15OQ81BFvHTgO/bSU/5rqcEhmynn+/0QbXZlvsIhn5Wn5Da/TL7GMfGUP9Sg+gjgusDb5ld5z9
QhBTwoU6WPPPYz2pV+O7AsrMFB8oMFHPZMNWUm3GkDLEYi2XH6g/ibwcbHkre0VV3Fbpf+E8Fd4F
LffHv9XwTjgyANBnu8qD0DqHIvyR/N5mTlTcksfbEgmasitA3eV+fwrhjiFBPEjWnWi+7hpJn8pD
W9xuEc3Hus7lh5nxiHVdDurEA9fH6ccqH8g8h30NgRkrkVWYQziHD15loFFrTmIE+6XKDeTeJ/R0
UnvUp3o11hZuVEe5enVXSSJmHx8lzsSUBuuON7HMOyeBxp+GbQUhCKNQ1CMN5dfeoi0sDA/Ir7uh
RrZbOgeGbUcdz/+mlIW0EBpVn0QEQS+0wS1QydFl+kHLLvEY7/lPwlpVpXp4R5xpg/Rj6eCLxG1G
7nm9cjR0r3Tb6zeiHG4AxVPJ1BVHT5l87z33J/zLnQVZkQ0etiJPN7/I5hCewCVmw+1AdMTOnmny
oKcfcO2XqArsx54UHC2n/mIJh7ZEINmdvhllxfiUOmzjUWNc/NGNJKvlBov4oLqcAOgNc0YJBdYF
W5+s053A/QEtfedHhEWHhcvWlixjkh3kkPEK8oYf67oxaRcrXmDI9RtZoUTONjcrDsTomO6vXM9+
TCxE8tHMiSRd5HPIRtqOXCzA2QMA2IazbjkqgzTb7MUWdupkWlOFhKzXQPCF0vdI51u1Jj4bM2/y
cSOftIg3pfqOtIwA+o/KwBntzrwcuFYRrSQeyQucLfmcrMx4aquMw4+kWv73yZhH+aETE+Yzxpj8
xEe+ZJzrR33i2DTu1LlE2qnrh9gJPbeDiVzCSc6vyd08T5r3AS/yaEF8QVrGaYBpCDpDABFjvRrD
4AkIJyKgn63a6KUHMcA7+LAxzkxa6dGEKn5lw4/3b3UkgimFgsTn9Fss46rGHHFsE/aiH5wAyABp
EGQLj/TxpmwVVHDZ3D1Tf686eJ+5b5NxLmDEyuJ0k8QZ3meyOUe4lqXmon0wF2dLMGTiNL9EJHUv
eKgQCvNq41XDYZ3nEBaz1kWgddp9psJ+Js2YpkgDE3w78gW+nBg5FUqaXR6uqsrUXN+wCWoOuzsp
EQeJuXUb1d8RsaYa4k0aLafa8tMhRpr6lWOUfs7SlaYn89PBzuh7cRs4cJqCivb9aK6QB5fj7jcf
ubnbPYvZ++6GXtKTFwLajay9FLgShV6S55MTljfTD5WbbD8c4ZHc32WeBzjFKQdSjVVY1rhfYP64
VjYyAcp4U2JDGydMl0lpsOAW2uiQ1Nt82lb1r7TUAlLPT0bwi7Fu53+iUBEHBcxc4I0TCAWS3ogz
5NHd04mE88RDAZp+Kpcr6UwmmqRQgqt1MphQ9LJ52f0CnOvVZlSx7zR09Roh/2tUDQ8xadQjc9k7
3okqSFIrpcQ6NaE88NAVjav1mAaHWxzFZkNW9Gd++wSi8DOKQkBR6Cz1yO3fbO6bqm2i4oCqnvna
VvOSB24DWHTaMjlSDVI7EDvjyJUr1eXsoZekrPstxIF8sFwZdBv6SCedt35xFsn0IaTS0GIh9Kop
le5njnH0/wQNCwhfcHcKptYq+d5GfTD0XbdJwRm90bsocAX6EiO0F7MK4NY1JMzgezPfE3szD1Ta
J1gzAP/e5ZOA1utGwmXTDW9+S9bM6pdan0SVwWDI2iiYrU2Q4SRTpysI5jWCmIBiNBEZrCf6bvS2
ZQ5eO3mtFqqwtnCWoRSGLxXrTbR9wq2bJ3R6ZZke4OxVYer8lOlSCseOD9zKrSD3/UEvPqbLNsTP
CW/z9BHpTLL3lfGG69ccDZgBGmou27+WydZAemk0RJanEm0moF+KYM2upWmSElDViMIycX57tn5C
0dJYZWRb4l8oz3lGlxnPmNVE70vyv3g50DgOH6B2YEISuBsUXrpCLEJ0UQYLgsXyI8pkH5C61a0J
W5C9X6CQPnXSpheE1vzWoyQBvci4cZd850Mi1kbxenZVi88sLkFynqkHppRJ4CEKw8V5dt1g1lr5
ljNxMQdqscVGl3XJWdhYwGZqUt+YjfKTMtJH7QFeiZJlQrgOojyp9SIKzAXftzClPRSs+E17zYoz
ivFG7jiFssGzwSAO5KSAcAnFwc5uQ+2yORCDLBvBO+FNzXzBCSZerlSWUA9d9I1FT7AIyc+mwkU+
pzJ6wFjpktRX2VOedT+qqemSSsypVZxZwkigP2kaDrcwEdpPZoVpEw+ec36QAoX1q1D1tu/J0hAZ
42LKFziqGpkAPSHa2YD/3knLbPZmv47UFcj67mWaquo94aXIRM7Ro2n2CY1qR+BpxS92c5yoJhI4
B9T20az+QfQ4Icdd5+1kaZMzpuQtJE0ruQA7ib/ib6LjS9NSf2qfSUHakP8z/Jmq/+4zFSt+1Rff
IcjLUj0u43d9RmPrGBufYCps4ggNM9O4N/5V7kfwSXUgQSO9DWIUOZUxHfecLAxQKyVN9kRIvij9
wN86GVtJIWtVCsALvaT8AyyxkVkPlfroymQauq7ghQzq6hUAmI3/nK+HXonCrrb4j/XJDiUgXzIR
kZDdUNBLf7R6ctBjY11MVoBmwadAaqOFD3dwGPZMraZ3TTAK6dw8pQl75BWg02rsPoV8ra5Fq2DA
RJ4/QK77y++UzvawqeL7wYoLNdrRu44dJSF+y0cpFh/1XUUUVkbSLj+3Iutuzsp+B5iwr3NgBOp+
vHB7H4ia3X4yi2KZZirjjqGxE0pMkF4TkxeGkEROgZhMPsnyaWaWZkFD9cMeoXTeZJkfGY7RFne2
jiKvjRC09fWnJyKTRynr2u3wjw7ZQCMEYRu+QomP76t4AYq3YajSGlcXORP/02TPQH3l/aTUkUoT
c84RNZB/rGvaxLwa+wIPLQOPVBhwZzE6k1pGL9jiRCPwDD1zY3dWkNSeUlrelWZaWEAD4qQ1lBle
kdD3I8OcZKq8mL7rDZ1oMF2PzEPCtt8xPIJhgsAdcwg/YzmKEPflllvxu+NlWJ2YBVz8XZGEUd84
u1EuQNxLV+lr/0+0Fmbq43cEF4t7KhwzX8lq9dRhh9cN8nDOaPoVxP9wOR52KMNvJKoitkHp0s73
OR3KB1Joi2B8/s6rGs8xX3/qFqLP/bHezPLSsTZk3ChYH3WzimSeT6gQ/Hbvtu/rJT8fyyea0UKw
mRhGOep5q+IF4xEEDV+emXVHaGKpLlYCBOCKYGKtTTU1HZxSqX3lYkD/J8tJ6rEU83EMlqVcoJdP
+GgcQegbxO7HL0qCe2rb01RKy6ng9fcoYfV+m/U+GzzZ0QgdNe/2/6dWGSWtDKRR/JQws7jGJkTo
fisgY5AVgxMfzuDZfApUcJrK9zSvnzS19w6wtUvTFwJdBbUpMpv/l/+62Nx2cCBZJvfNkfFHhZX1
ohKjNGoEHDGW6DFoYAeIYY49TuY2LIdCK9Y9ddSJiVaEd7vba+LiWNjRgYog41trXtzkukW2AY60
HcGugudCZjkIDSwy0oeupI2TBZc2WbOL9Fz1pVl0so63KRzUJM+I8JdmTBG/kP1Nj/YBZuY8eZzC
X1a+W8K7IEz9uBkprIGGu6hR+fO7SBUuR9cJL/kUKwxFBWQeLdCnnTUKmTXl3QEddamGraej28Yn
/xWr1F5w5rkXGWg0Y+wE5x/6UKddR0lyirVEoI38pmEfvIYKGTmL9bzzAsgRuEgWtIEamDpuxF3j
o3ep8o5ofkVj98SEvROHfDtwq+YfvuXWT/W+pSzbMZPDWAp+ttcD3Rn8QEcjw8RSZFnQ2S0yK0yh
ivBcVY6Si9DbJAoHzuX7OilKlAhy413/0+vf1PF+b3ty2XhaMnoepxlVG+Yzhs4E8l1c3iPVZOP5
rhzeDjZKJoxJhdvcBGXxIHVwISxsEef4ktygW6If/VA7hN1pSzZazCqnFlLE/bX/kiAGtnY1T0qL
NHGs6r6JIWPUObl/kvJ1JpfaWZ6AiEuGzgXYW1Zk5GHd/Pt9AIqRZnNNx63fDEIi2SWDiM+DxahE
HkzhbL81y/mlBH8o/8G3Pz6eOePcfZONkV7jomVE22F3Hgelkj2+bgFK9OdLulsfcn5jrIcY0LMl
E3MHIfF/cPFSPmYB6mfXoGqjYGUZEFs3NsQAH/JBXSVn/lwPtD7bXy0Do2UduPaZQ0nLIcNz4qb3
vfRWzVe6FzO+V+EtIrTwNFfBYpbHzzI4TQKdmpQxEZJ/lRAbtTbYxTh+uNWz9dQ8fq6GcHKRIGZ9
I+umxgTzcCA/8/nm1YGSv61HZ9dMpWudV/OMVVC6rGqYyrdEl0Gqi7Ko+y7yIOBtatyRLxYcJG6P
og96ZYT6WuTKIyiKBKBLzOriGbu+ZAsFxfY3536i3KuSbg0ES9dQHj02xElf8NYdSXnN4b9E4jST
B7gMvQbeWoaMDe+LHOT3KEgVQw3N5K3ILT8JeEhxdKBalNVjYMge3bvlvInKZMAGfHy2jHOCFBgn
3TsGP8Fy50v8uGj5kbKqWhbjjL54pye6mvBr/Vy5tGVobGTYYUR7wDLwmYE+vQj0ELikVbVRojxE
jB5xInnM7CJTyujw9iOQg+TTPwhowuTC/OXiqYlSYzOkunB3c8kLPvVm6iE8n/oW+OsJrYFysfX7
l+Pcz31YXn7nREBQiYPsMT2D0LTvMHaHrg+f9mUDynxRT8veBTU0GSoUHOxiMf2OgnfLDcBd9mJh
y9wQCqHdB1NwNjMG1ztOLFnYXn2Rw9qDkU99hgx4k4bkt8gnDu/7WkGeAlZpiK/IyXh8VodoOG9h
cJw8mYGtwUzjuwExUmITKvyOzUclYuQ3/BJzEBO86DeSbzDhBFP6N0Cgblbh5rBo5JV/GKOhGxxL
y9LxnUmYF1Syqukr5nArh27R4yT4fT5c0Wd6yHtZHFMljrGieqiFV0H4uIst1ypISMe8PR/6goKO
HqzJdzF/FQ8rPN6Gpb/+7/mkzLg6BbPFZkJ4J2xg6EvxxSYouLY1nqbw/korPrF46wyFqL/jTDVt
HNhD3QwJh50Kr7CuqlUH9c3KxR/V0pXO7smvBIBO8Q+4ZQH0ovWZOcldUS+yWMA/ZVND/y9IV1X/
1kyeNT8igERjy6jkHmWOy97HCqEA6d++CVG1kPZzLT5AdEguP1e6LFDdzxjj8dOzdcSAMC3pOtRw
CXdIW8fKfa2YL4w9lBp31tHl6L0ZQ6Aq2Go8HNPh6NR+kx0kvpaVoOptsQO560vrJ+hq/PUIuCr9
WwJxG440blAFtCJjI6qzwdWPm3+gPrGA44jCNnG6PWLFThS0gcbCoLePE5+CQMfEDgTgT00vopRL
ALGbrOtwdT6JDCyAGsVAtjHye52vKbxYvxtml9qGMaHs/mEwZoMpzm5NrlwEwxCbLFKFZDQmaZVY
7iL2ZPNpuhVPtIH2Adhs8nazHT7Uw/getPRv8yzFBkOVSEwiBObafwRukHHIKFVr8AONV1IJLcHV
Wlswcl+y7iTuahqorVPcDXwCpnNfFJEtmuqQu2TS50pBUevzFBeFb+YOncXsZ76iu0/L6Dspi5BF
rESCeI6aSOno7ZtzfJNB3drPmklM4N1K3cZpLoFc2KGMbM9waXtKLdqRwnrGO+ZJKk1EynxHcP14
Ha0edGzuNd0O10R/uDddGu3IMSLLDtX4f+TkUwOthm0KteyJji25xslh3zKHnIeMEcIZGUn0OZ6a
gAiOwmjmR4ryeynouYrtghPAjGXgjYABdxYxnNcJ84p59XiErxdCMSZ4uyqbTo/lFm1JT+hnww/t
vusLX2KAzbiAkOz6Hs6bTyJE2ziILoJbljCZ/691eQnuUhQhGBR44S9gLkzLEv7hDR5mu5dh+dDp
Vx09DEXR6TrZPr3dnNR7/9tA8P+Yw8by30EA6b6G5Wn1FxCB0vgO4yvsKMceM9U9SzGa5rbUE58F
6wAM3zGvt3UvqqaWQYdqTrz9crz2BEfTwIAFc0zBfJiCNc5g3prHgIH9CVgMWymYgaVPX5AFD8JR
ZTo+z6G/YZsjDQour0EzoJ9LoctWLmSrNZCnyL8IzsrdG+koMc0OhHei/zJfSPmH7Y1lrRZRkgCu
Bjep6vsUk4yA92uxsyx54g4IMoYcTp8ueet5eJyfEzQ7ZH2SVTcwZp35US5+SYzFuk2V8FnU1XYx
YzpmdV8wixLnJsNpRg8Uso0/T3i3y9xs+I2rTw5P8Ugrqn6yg7NxK7KatSR0ub9KmLFisXkHagVv
maejqkXwwaeY5ZHp54s6UJBcipjq46nuhwkWTm3Wpa4fhMCjMVP3m3vruIuIB7I6IM4HIc3WJC7K
ajmx1TFFJKUMq11rZG16/1gcr9kHXKSnX8EGrSJvK7lYUfkIls6DbPyMxIY77XcIDZgTP0/+6wco
TvPssfliInnTZt2VY0cFcL+gjn6oXi62HIEIrxl1a9RfQ3C57SyEgmYu6xFfYv6DYku6IXtpbO1A
AyJCzyoxi+PnLiebEtnWo7jvXnGZZSZU2JJxmXzXSy9f0yLzwtMdYSoVLJK209zCw37NLk8OSmsM
6nl7tvxYvwRaBg0T5un/hR3Mdqcx6kbW7LDGRRfzEEAOltu0P04W+KghWxMyFX2VOkoQHvyBsueo
X+3L3RSg4W42FTUcYR8iFWylaVXW1BCgwHH/8w4TIY3go+M5BIO5/Eu5Ye7oqf/osf4L0l3K1XB6
HOWveOWNV2Jy8rLU0/NpMIp8Y2IFL5G7YnZmShcCl4JaQyrQdTU98rdZmtU3704ya4Zn+CZHHQCS
gdhcRvUZlmc7o3gCT50pSguZIhrJy/BXzP4fmGugMOpJdzm2O86VO0FbO8r4nN44ylVKJIxzIFf7
sDDct2FJ4XFqMd1TkYkd40wxbbGi2lBMKsCt8sK4FKRoV80j209eveJ4NyMz5+meFknndvO322YM
pIXI7jlb2N2x5jdokG9hgflMFArWLjsZQc0XcGJC4OoIm4uM1lmfZuGiHz1TpdyiTqAUlzZVHk5y
3UC055Mu25djWDhAYhmDqx3SV9xJq+vRykub6pfL/yGojxRAlgG7+hjWeRgejQClifBWahzmv7AK
LLqjejNqYma1Ew4CR9SlYQe8l3PLp84yUFpql7Y4zrNDObLrf1Q3uOxUTbGyQLfFZWSFBVy5UrxJ
UKYU6XmvyhJzG4ZWTlZFf7AKrLUAAFt72jDKiJniJoFvb/WsGicq0XnHY6tezLV0S75te6dtmqLJ
BzsT72PwagH7jc3zQ2Hi2O37oFypkUmK1dXgfUoW5hG4CAYttu81H4LI18zkU5gwqnhp9ZlbVTr3
BnmVb6KS4angxndlmkV1Jb/I+S3BQQH2u6DtzO4pG+4hIRm6ewx2kcI1XHIkXAQ+E9/eiXThZs70
7TZxGM/OU9mzOYvz5swJsqSANq+uLdURXDbt9lgZZtbkJIamodGXWnAVjqRBEHkjpKEJDzX3XIQG
ZCF+zrIOCVmLOFnzKeVsEczS7WKQdg1GO0b8L7AL4PE8ABDT97VpgO7OHgdieU7dJh7fESafNgdN
R0SlKAsuSDndYbiZ9BopN9P64eOX5GpCN8T1y//u8hr7DO4kci+WLh+e+pSqYIxowhPyv/cZcKcF
cbvUIIsIxJpC/DnjKPkOUkXpDrCoLdTfGKC/s16wnrMjVxmE/5sje81cD8OI9gzNpnb/JIzHW9+u
ueOYUsy1gL67cQ0CpT/gMu9fHEECEQJXVbJgThGDLmV2JXHbT0qX1uZXhc/kk6p4/P6EkzvcLeO1
vnlxSY2Bx3XGCoshj5lUveoBjnTsegCieaZXAjLMF66lqWHaM/f5Bs5sIyRa5b3xirTzL4brpfF/
9c0J1/r16bavLImvImZnA0hL42DkJtbZdd7z6HqWE71QTdfwC7BX+ehWYS8rPpIGp/B0tgsORZen
2apKBVMAM0b+LwDuh/D2IKrIkd6LVoY8EKuv4o9Yq2EHgxgsob1XPLiB8UHQLFYosIoD3MsthUCp
yr7rWHUK3xUQv8hnTJEcg+bX6/b7m1ru575yEJDGHqf/GM0hHpK+cOeL50RUmvRW/tPqaPiVWClO
hXsl/iTLQfOFWrOP8I05/R6lz3qSii70XYe+vbKUYM8qPXmj3hDioFTXGR2cy83huUU/6Mxxrx2l
qer3mYFcbwmac5/3Xa8RHDrOI9/rfRqIWcVoVIgfVdIdGW8a9dQhbE8iIBobp9h0+hjAvDRbnkGp
IX+asdggWtMedHd2zZoJa+R91eYl3ubRGDFPkSWKkIXbBTiEE5L0wdcxSFffiKhhATD9ISgELYIY
ADsXxvMauWALA3rzRntUtlKZZw8TSXw68XkHxHZIwjN3oq0vLtsjeFIWyzwT80QPcHTiv7vNMqHh
hD8o7X1Q7ukNcKR2nJ6Ygsq+ijSBkQFMSlDHeLMSSDTE/01JVMCjkDxvsVKQKW/X0Rv8248nvFE2
EdU3DUIshxgUNvV6nMMzbAEM3j35KFZWtbk8czFdsyK5J8MdquUxa2OwgP1UCW2gdZPedAC3DgA2
g+lJ64o8A/WB8TH5a8fwvXmosOr39kknIwdA5lsL8d9DESryzgHlzHTsWLhQf4ho6Gp4RRa23Wpb
YMd5hikRZLzc7R0s1Kj/EsswKKXBhr7qlCacIQwX/mT2R1S3MFdvFtld24tOWvoG+Wq/sbD8TXxv
7QZWR8/N8umFzcvhJcRKOuSMOBOcWWaGDgnCdXlYxd7qCZAQ/sZwJWNIaP7cl3brdpNqpKZIFFOS
tSX6rr6FFNiG9KvjcpOudG+sRmD1ha/8uFKX0DPW2sGY6H2Zk/fW37n4VYITXXM2oEbux0IvXPB5
unH5ryLbRKXnlaGP81tcaNaqwVqBmiDKmlNsQVsu0rMrNoa59wuRE5NzJHVVWllw2TAetzZ7zUu3
h1P8h0P/vN4lwZ0nvQhXFFqOPbYPNM9Y1+6ILIO21u7RO99HdyjYrXzfl53JQc66JIRcnWuUNnq2
Ry/GNhbTFI0RIfelC7hPMjoIAyE8tzi21IMVEFlsExfpqGFdnGIziVKjwCl3ddsz/B93JNIzdjhT
rKixwHSx8XonLYq0yQXATI+JTd9GN1SjxLsLDvMBNa4wjUG3AljSCIpcIpj2hmrtlTQi5mYwgz7o
ZUCbFQ3G3P4LXOPoXbf8of7r+y68F2yY36al3ekgjcEh0/5YQ5smu+G6UiG7Pd82XMn8A3g65oW8
sgkxcn/SvpiOTWeHRyAgmxPtMHrGkWr1Ep9eHzxANXIplY5DkdO54enfodHA3dPf+I3UgWhyxuH4
a8YOweqjVBrMFCgNst3gcvBK76yV9SQ/bS0rfleS2IE57Gr3/9phlzh0gv11tzS4oFq3uzi6ZthR
5QKRFZsAMKgyvTzlhsMBNNDeQ/IkSV8GvX37uIrob8NHKxgOik67IdcLzIbhw1VS1EWus0YoKRCx
Ra+uB93WvuM2bkbv/CCHm3p+pOxDdJyjpIjznPCO1B8YbtHlsBU8BciOk185KbWnwtVWvRFG9gy+
kmMjHZEC14Wx/c9tyMh7OII7JLDPtZOahIvHT/j8gMCIsNJtARQxgPGf1EDf85IQjTkrQvzgbg4V
x/QGKCYOAnJZ506rBLUmHQCVR/AT6rXWr2fTA5EyqLLzYy6565J4y36DJ1uvuUw6hH9xIMFIZNHb
eSEtK0laKjdQjjKkjhs9F2TwoCyZuwI05GtmoTFwVlSBQdlCYVtofkHK++I7KD7cR3LE0++4xSFU
9vQhUDdpX/6Gz/08KeomSSroll5t2/2yvX0xwCYJTlbgtXqfHP69UJs+dNdaAMOp3QEeq60YxnI9
kCeCuzl/mW1FVPi4BRUPMm7NyaKqRLK94DBYEkTW7O8XJWU7vBZl6H5hLnRYsewPD40UwuIyY01o
Rf6kedXWGoXwky2bTzxycch0uqKnKJXMnB9HWfd8xDvh0NBvmv4mM5c+LvbAQuhw8lWkbjRcBDly
/Ak9LK4+42Nja5JvFqwDK9BJ50xB5PVxpO5+KYogTX93OoXU1i4sTYg0vVGj5Orlf1gXuVEebfwd
PKbkjaTYLBuCzag9BqYzOOZw64sCqEHK4vX5sXS8Q16MhRFtOKOdgFGfxXqlppoxnf8FwczUfXOL
RD0Nr2SW7P1VMFf7FtauM83Od6I6OOD69eI0JgICHFVrKoiCwlUrLjWb3eRYfHTmENQxp4n76uev
B8+ODNY7m8WMwoOx48y0VHawD94EYJxobYY49iCdHAaWxJpQLBiJO1wTlJaHmQs6D/TpPEPSx3NT
UXmGvPNajiNx95mCXLtBo2l6Skg0qdq+CeENGuxn8ZkDREsbvqIM8G6G/LapU3qppwzjQ16voQjz
C6kc3VY505MclLbXcrFkh9GEmbkt7ck5s/AWQUw8d2I8NdaDJUJEi+u6tpZk+i2B5nj69tNlhbLR
33jBalniSHUrpZ92EOCLhXYe/wO6iLNQ5NmI2zZuALw5sM6xNjjz9bIUPi9+eSCTn6oBVFfDTITc
GNfLxCIR+jKV2DXTW2Cz/4mqKCYaro7Gj69ojG+LQMKtwEss/5Cgm4BAXGFYiI/bAl8mx1mN2bCY
jVg5L/6fCP8NzDS9SOS75njXWS/sbmIRmuhhkNcnqJijQDywjU5F+EAcZPlhdfVJoezDn9G/iMZm
Tr7F7q+R5YUgxca03XM7o4elAryAPSkuJ78xD9YdE23eVMeHgmYGvf0i0Mw2yntTgH5P6PJlkwNN
Y+HKpesggd4/sc9RRlWe0PNnnjR4ysE//ZWMW0bSgTyGsWQEmqnojoYDT0MGHTVckCxb7Q5sQLzi
amWPyjZl7x6XKkrduMN5mHaBd1VsJndDzwGIshYRSpiI4u7XK4EuI8CvbVFFuJUD5J6dl6A0yYVH
LM7OWWVluiQQ1sq6V6KK4gGredUuEtcRheyRO4SJD9I4+u/lpv3oDQEjAWyh9cl2w7mgV4gOpXsj
i8TTQCPuRu5UnwH8WYjfwXqBLj+sz/F556i3y8tSnS6Fu617W21b5Wb1n0E0bE1ao0GXa8QlNGMp
ziw8TTlLT4dFZEHF2+JjOAyeTSzt8Z25Tb3Nt2pK6c8YOS5v8FNuXn6TmxO17eUwGbYsLGAimymS
Tr+WSN2u+12ElS2g6Ax73n6vTLb9vSKwj5C85q92QzNNIQbOih3Q6ihUD4/7miKUtsrzBC9Uwfol
L/2LWIbXYybosGCrnAFOdPrC8BF6IQH9PLZNLtB39I710hVjunt6OLAEaAee1BhxmCfVXOI83FSE
sAGcWOXV92/h2VVLxQvIEzpbfBFMnlQeokqK3yGrp8g/6EYuj9dRi6iVz8cIe3vzGdUeN9wEUK0R
QkEFUQgaCrD71GIsp0FNdondH6MY6WXFYatwGhNgLfZn8fPgxnEzUY8JN1bk2J/P2epItwRGzZMA
QST+5/xmW1/dqxjT2yq7IJZu7t0ZGdWlDS7+Lv24NcEVRdql1+4VbSpE+ispXDRcZkesczFBVgSa
oTs/SSK23pZ9D9ZKLppgb83u3hi62Yr867nVX61ZYk45Pcz9JOfF6PgB6q8aW33a+4erdm0AOcPb
6hUHi3GlJUnFE5gBLIdmRU2vKmDtXm2fJsH4wJuhxYDEexhDDAEuHj/fz2b4EhAxNeFZymUj26Hf
zT0HTLrTyLTubH7LGF8wZkthi+3GTf+9eBdDNzim+MP0y8ZZ9v5/LkbxzBt3Cud5v2ZXw4X87X/d
0PIb96HVxOwlaLqQSodZJB3+eRM77MPwcqC5Xf4700A03hlsM0E6fKlwbhJySP4V/tfdgBSfgaSw
b08QYTbUUID7OzvGRBF4YMRxpr3DH2jc+Tvt6q9RT+nh1D5KgGC/BxrgCZnpqAPuQ5Ms+YG0vslY
/v3Idx3AAkYdqzQp8M5DKz3iaDFDL5aBob+6cwg+/+evvvhr9pj9K61vD+b8TDpn0Lg7shY44xEx
24VdHV+9/mPG2HcW5kWLCvA7EQ0JsTvJtE1zKron8cHi4DkoO9ndJaYsCQAAaOBQSugAX9aaJGQA
r+94e6CqOCwqA5yDwwB2Z3yuSPZLF8mg604tYOk8gPfL868G7Igd952rsTPUXZQNXt2MEZy2hB/z
fZBta44xq0uMK2pK3pzgZ7RNhE+Y1QdNyaCb5vjlufIXlZTobAFQdRz51Fuee/unZGG256M13r9r
ar3uoMf7ehlpBa/QvFbp/sW6fHqvkkTnvuXJ8Pq4Es5j4ib1aU5yIpxZMWfXCO3+564zcG9pr56D
qG54MUfKuSLGjEnbL/6O4ir760Rhr5upfqGePpPRATGMhCV45lnyTSxdXkVBT9aJBMHBQF+j4fyr
3w8KisR3Xn+lhVzW8jZNY5CutN7EgUCaeJb3lbaVr80QmxNidugKsLzYaIoC51XfLwNUqjcZ0Fcn
KWSZ+JVHhQj1BCHwlY6V3qs+fUPqsOBh1maMQlYYGJjaJOdszHHkMIRiZhqj7kVKR4BIC2YZGjbF
/gLLIBk7pXAWebR35WKGEk3YAaJ1QaVTPgczCWTfbZ0LGecTJUGjPH2Ir75oIe6VjtVhU6Kiy11x
NDgyUvJQX+3Q2B990/X2a4vmFqFLlybJN35idiKfwI8+3h94pzUjEUAe5hTxxhb7eZIAD5gwqRtd
Fbh0Xgnzu/l5kElC7LdhIy0m3XzG9EVgOZcv7AYW2BrqrpFW+JAinpFbD/9xJhgmC1HhXe0KzWWH
ieQjuMMsckCVEDa5jzhQ1zs/3KvunXJOqfQ/5Gh5wN0F9jJbz9m1laldSG9VztxOKZkWFH0qAGtM
KHcCc5Eg9yPnfRxluHjcIzcJzPU7kyYFBwPzbgAECAvPfHjLjudwT/fpcP3IrpTmnG/9i0JjIzIv
GMxctTGOLCnYHgbp4bx4HBBPUOY4p5QFob5Z1ukfpJEm94tWmH7TYx4bNQfx//YjY0KFLHULh2K0
9zzS0RkiVelbUl+0gElw7VsIgRB9f7LMZhyy3cJqF0Rw//9IcsVoiOq2sKuO0NraSYdidkVknIyV
a+BNa4CSQktli0EWnRncbmrQQ0sSuZGNCn8hGjQ3CYj/Bj6K+e//gAxkfDmrkqtxD5ozD8CHjr2y
lJG17nxBxPv/51zm8s0I9EKARbR6vsgvaaPY3nUvTHZiTsCVBHoNkbTo86DBJg8mjHJJfQoaqyAI
gyNjybkJxYn3myNIgiLVnyWjh3TneDTMJaxjrMbiXNB0wHx/FiWlJuZSE6AD5CoDs7+Ei2vRFK7S
im3nRQR4mtRA9gCw7A6bu924It5NdHkbIHsKsxD11c7V70GleQu4BKJZ1xoywyKBHXjpo4YNWCUf
sciw21vs3LpjvCsLdKVRDH5gxW785rs+9JP7mykwzdcM1ubJTs17prOZs9vhxx/7waFFAXdbQxct
zDBejn/DU8SU1Q2TK5DF7YFdBvSl6D5e1/QhI+TGURG3ed39X73ZDhFRZey50A+ATr2kd6GJ5q4M
EKNjfDzEgaCAoScQT5wCcy3vZotn+x6MKlDGVIedGZsu2RBjNyQ3rf2Jk3Pn6+bKOYtazze2f3nC
PjfyAlMYab0WcB5ckQgZ302gykba06tt58thI7in67S6SRerlL9fAX/aGlz+Bz0CpfhehzIKUwBL
XEe6e4N6mJB4QACun+VLotDH8ZnTKuasHgohLKh9qdj0HTKMGJyetE7CCyje3vHQVrNOROUj2oKC
nFckDYotjF/yavesi2Zec+WfkZ8BfQEQLrVUqABAayNbpDuZZR8njPQrj62WfTTnO5gwf130duz+
2zFoiBhoVIMAa5cN7Ilf3nExjt8wdouorqQ5F0qjIjX/No1Bf7vVV6kh9HwWw6YsXkkmPOMYu4hR
pIfKSKriGvUuOhUBdplcY5fdTihmcoFtJXEuSNBRHBjn2WsIxP9Q999gZdZpDDC1DvARwGY2DFB9
tJnOrrPEGdpe7V8v/T374ewHiVYBpG0YQ927OiYOfd/yeLXavjPmg2iJVlkiFK1F6yGUgDJNapEB
BBFiVclG6KUG9+gh3Lkcg66aFW1457aSRduQWI0g50qcyNug5I1xvWqlUCpz3gUaDOelB0zbj1Ws
hn3SRH7g3XtY03gvHUjqsbE8czC6UZcBSxK6uAVGuBzvzLO/SyYMpPaoKoWA0yIzpwQKCm0I+Nv3
SfY+W+kHC5K/1W/eV9A5q3GlCDvG7fTqwgd75cDKMH1iR6Z6u5pTdmwcFU072vg8UQ416tqQWbtx
4eLnZj0fLonCpTnBjRf/35BXtPSQyhnBX1xshVieqjyN6fjGWcFpb2KNCTbcvAlHj9edvEVKQa0I
Ma/v32xbjxpKLUsDNlzHjiGPU8tZ+645yko7+d/NSKqwzTzKKOkbH3aIlRkcvztZ12aMHfsFMAz9
hoYYblzyzs+6Sc8DW8NrTvty70rfP4rfROBuydTuDlzsXakJwO3PRYRp806FOMjlpYUtrmvQdl2v
vG4M987ib3lZnLEiq7AqUCSjXsBtShsRaklrww8/9OQ6mPBVhYA5t9jTD6EnAgjhjikt0ZZsY4sz
1+wJ95HzU7bBjcAQymSOBgox0ISuHHIjWgWNYUSasa13wjFUBA9nAmgr+G11I0KSpNc0vF2U15/L
irCPZbZ2XqsBllamha5eXHQ7ichhUZeQ4mh7zr4qNgiSR3fNnypjdUwHAQqlqfeIjcWB8pkEJXjX
Je7INmpvNd7XodHwm5AlF2ehRqqOTuxfWRmfW5UcutEqsIsFGps4EyCmbgmamwxtEwxBUPsJCjbI
li7pex7crYQTW5QizTuApU7sXGMMPWbJKKVTRs6IVz7iYqQnz4+DHaDcM6T4I1DjVwyw5KiqzINP
dwHpsiZF5aKCBl2tFHBf2UJx0xKitk547xqCKyIvzAfV51foAD25zZXhRHXaDjPnZUYk6gZymo2o
SXzSDCyygfL4ja/eHe6IfAJVhtFemhzAyePFQ+a7j0n2BB9S9xfinqvKTPQbq3QbTrMuJ2rGDrmy
24tQOAFoo0ZluGligeb4Szh/hG0HYWhESFQSvwxpV974zHYEicaPZbs8+ZSHGsqZLTS6mWu//hPB
SILbj1U3UVQs7qNi5URaV0fQNbapYHUI/BM9nLcB2cj4e0HrogZgqSkPqvpQGQgh1khNvxPl+nut
6Z5BCVS4eincXFbokdw3/QN9esTyk0GzyJxxsyv36FNVCEmMsa3NRXaiyxM/S5tAVpKFVL42ngtD
6VRsXcJT6fqPo7ZUtQ4irMg44v7EkHdknAm4MfVkCC0yCHznND1s+x/6tJGtjCLiZO1mZUeApQmI
Fx33keqCth1jUvyXFHGZDknRmhXkU+ad++NBxiyT25swDfMiKzZWdBHZdVrzZkCF9r4R/Ka3M/nF
oiKXMZq+gQZblIsI9Ahd1TizVAjZst5f2/B6mZfDkaL/yOmM8Nti/nNOAGqC18ZRcQ4G4JyJ8Zxs
ZjkGpe38fma8XHmFvLcmPsVyalqVqq5MaX3Sc0TE8U1CJgTYwfnCim6RbZ9303pL/sGE8j70fezN
r6WZDAhXIajk6sNlTIvcXzo6jyXTMpk+65/2+Or5MXiZaUw1FgXKkNJ4t2WJl5ye+UCiKHNjIjrO
fDGOUg4PVlIwl2nEj/bfHGJGuw0nlJA5Yw0lZ7lDB3WiQSHv3CNEktcMwnuLPNbUsKxuvx/OPSXL
K38TOPPKwXKqDbrEgLFVjahTzLUDRtsrLn5qUveruI1jTMx2+mMRwb8HW3X/bmAlJ9hzbNEdkjZZ
CUia2s2X7RXlarkghK2E2BOyHi24A6lM3EoA6A+izDGrXpc4uJvq1JYallesuaZcybx3ZFBXY/5o
cbxLGld235IqPwguPsNLFDKUXx+Sc+uXhv9YS5XP5dw1SYJ0XMDLM0sHyxdrGN0xjBeEboE8xxy6
eSG85QvWvdDL7DMNZHD1mCc6X2RdWmyjkr627VQhEIlknqaUVqA7JubBqErnBz+RFWutu2NvHDPa
K8oG2neI8uBtScaKuZjFxR1uTzCT8P7OPUoUJJw9MVeunjCr130JKjQyeMtfXwGseFSCzrzGKbZD
BIAi5I72GKJ7VYjyh9XwtCveTsIQQ/2pn3d3sX8/Js0ozYDMlGxb/vlFS1LYt+crlafki0VL+Ksp
LV0Gv5rdxQte1NO06u1YEnQ4w5ACNodBpfzFpM3ioXezRrobtu3btkqqTwSiwsGjpvTVY8MhtgGt
bGbjilszuUlZP6zNsoD6z5ypmhz1gg91z9YvXjwOb9Bbc7VOStGrHI0+Eegr/CogRs1TV3kvxksr
3Y46XzD//vNOmJdS66hD+wIq1U5WnXer6vdrXLb8c+K261elqNZbOjiv23lRql2G4qvpjt+dvMZU
vMNwt+AW/z1hnbEwnBhyw6v5rYgbv7ZgDaLtAe2irkB0pJj8o/Bs2JkZ4c/BzgEG8fuCtLj/p698
y5aMleVB3/W0ShwvYlmQPbbt2mZEuTe5uLaXvk01f2AoffeLP2TlkGkGqnPjs2HrY/x0kfhpFOpI
ZD+INN+NwYuWLuo00u1g6I7Tk2HgnuhS455uEvvTI4+4YjQ4ivlEAEsvT7C2WK+2zlO3fO7GNTvm
u7+Z1N0IlN+g0gmCdBaI8QMM7Ij0ByVFYIPQyno766czpr2lvGSU4DnA4lSDjha/OPgxYhlqFMpV
fEJDbM1grJoiMDkZXXEMMbGvUo6WE4ohKdW2T6tzeiSkV6Zo2ythumuvoMhWRa2GlJCRqB9nZ8Jk
Fpix6WrBcMDK6QQclWMlePCDEXhDrlKtFNA1ieJ21N0I2BimQd92Sua5WcPzRzxV7fHWn6Kg6SLJ
GE0gsSDDVTsnUUN7RvAEhBHXmVtfrYUkT1OW0Butwu/A20CGT82co4l9IDpaQIvnmNajHS3KDA+P
+kfAq/JnMQJGK0RF837FfcJEasLYI9LTrSqawcePqmkyRaWRsV8zJCM28orhZiWSDrcjYnKsk0hN
meM14/AMz5BNy9iUyi3hbRw6BkQHjP9rXlUKJ21RMFSwlKOWP1SwjUwVVHUwUal929qS57FXRSwF
TL3YV3+WVucjhM08tG4ASHAKdKIiqTPkv6dgAZqJggoeIMvOSDdfiYzAXDLo/9RoHdMz1cbVGFpV
wnNEVXMwAtFlDdoFuQsLosPYxO0Tftu954YGRyLXScCCVM79kE1RXOxfg/EVdQXRp0ztx3eG6337
d7XFnXe69BKmVpBBbF7adFWJiPCw5R7c4LTujAtUbxxwXgvYwWDNzJaBJwzO3+oxWP0b4onyvu1F
1woXkG1qCsc79R8413a4sgjm5mp+G+GQndBR8cac2lNjfftzhMPekSP7NTyWheEOI4tWiUKf8kqM
sN5P+43PDCplApBDMwfsjjyDk9KLxaTjBC+5RpdrKzoQIwy1hZJOFHnmzniowXqxW+W4zYLGzH0q
yssgvxCxh4yyrdLem1N1btoQN/cPa0aQNW4vrgsbp56/2inAKD5DU5f1VseIkN3H7CAZpSjAiSgx
2D9bZeBRmhvBmdiyYuPY6ny7Aars5LUSLTjUmult4nwjBSNmHDdbVijA5ic4xxZlEq3G9XV2DqqG
nkNvgth1I+WIuw1rL2gIfyu3eO3mFJxH0ITVhrSPCgw+X9tUfxSGr9VcLMXTvCpGxQPlEnhQ6qzK
8tH5i3hVC5k+yOotrT0MYKyoBe64hHFJQMs24FB6RMlhWRvyExSR3mZQ5FzQA0/MW7Rpj4RMP5j1
m7NU651JPPt+sMpbZSAjC/q20pxce7SfAz1nDZcDuBpNE9hj1fG8xqn2JkFtVRGMMYhS1bFieCgb
NhwhC4hhTqopsxo52RWKlsqdqaJ9VoCI8GznIXiuQbD1ZEliFk7noslkPYJebeGLQs1TZbW8SIRm
wajo7r2OAbXZvW99voL2FEmM3f+kVsZym/O+XKhJttv+cpFI/IumnthrSufOQjTNJJoWqQpnlf6L
493n6ywM7NVSgIuSWgZuymu71dx6+NZV7AcSRN3R1CaOraccjITvbzdWda3fiVEVYXpZV8eY0bTT
rKdsydodbpQniw3elnlkohLOvhTn2mrzzs0uMaBimCxLnw7Ga2t52HdmvhmnS/6gEOyqq0LDuFHS
LLZMScmcMjEzNIXjwePYnrI5iqhyHkGvJjRD3oI0W+RfxEVat/HFko/WLkNCy8K5c/pXUL/tfW/m
SQGmiT8B+2ryrYIBHR7ah5Dy2HbAUnxd5p3zI/v/lsCyMIhzGLfzUC+cqx98jmDlGUVOg/R8gXDL
ZllBAkiOoiFubGKfaj1ABIpiN0xAM+Y+TjA71IjwiDxRhrP2wY4AzRR88d/o14YdZiE0W0SzU+d0
0Xkv//7zwc/B04lCJbp21cgSq/Cvz5l/ZoCy1T5w02lx8TA6uD8rTWTRqbVlF+wtEe5+UQ7pEs4G
1j69QKC8DDzOVeIAT9T8V+2n7pVXo56qQ4ppB+p47HSapefiwONgIwzPp4GK4BFH3YIlilrCV+/O
KbFQ+z08B6SdqVOcBF3YskQhjN0t1MB4Sm9sHrR5hpWm0XLOVVoCVGFr3bD7IY50PVW7n60JV0+j
L+qn/QvqG+XLrvL/ZDXur3g88RGn+5zZYyZEEtHAdzr2j2iQ0O9JbZ+c1RzP4tqEAWNCxqJlxZng
kyUqGW8vLRcyaX4nbCw4n/B/UZ6u0DpbVEhqZcZayoKOA8iB7PNHZhLbLLe3J0O7TCmTq+TjbKLR
EOkD6ECc4IZ5q6E+xZaYuLLEAqmjsQTEmd3M/jxpUxDxm1NTUCyrHvIp3ht4E+sPPg3AJR0D9fUF
hMuoE0zgu6vv1H1fmj2i3t+a1Gyr26oI4OQekm3W90nK8cabVRBUfkszLY2K7H44+8haqvuBIsoo
eGoF86iKiJXReA4nAWRcY7x9W3LDDtD+z7x+fSj+tWqOlFPCYA89gNhxr+b1yu0S4UQbuR8V+QxP
IfEMCsNSTExSs+/+hBJcklYEku/RwV6XszaRLY5sJr6cMu1mtRYKhEkQEyyR9PtGgG9CI2e2MF8F
CpGDL/HWEjrb7NUO7rmy6nt8nE5V/odUDs63YSB4tiEKsnERK0vFuAS5n9KGhyiNAVhFSsefuVpw
tD2gnYrx0ytbLOwMJCAf+pU0oWxgu97aD9peJMYDvWbv+iurOHC6hH7qWa138alReRWgOe6dSiLn
5ZxfRqKs/mkROpmmKQXYq3tUiRihRIEGF+A0DGkPHvpNiQDFhdotp+hQG97O7698wWa+2XVc0TlV
aDPa5y0BBIMe4xINcP4KxkF1zbropeoUTioBK30UMV4rckOOcXI6WncpXtGDx1T/eetQGDgySEpR
ZJwQE/GMLmRoVd39iy+Zx4XDXk+WtKBpLOemLFYpoprVWjHl93mQTQ0rjaz3zZ5xeBb1aluSnakI
oNlrCCdR+bUh17Yh+XIFpmemOw49RKKxe9WoA6kH8Zd9DxrdAc8iKRhpQu678Rn3GPQHwiptvX9d
K0AMU5g5heRwVNIHxbC5sQ9fdTbrW5UkLXbOOgTDLQ342qi24hqCA67xMf32CWegUgsbmZLW8qO6
1O6RW9hnEdDwyIqPPSMUtU8rSz5oe6ePAECBfC0vWmvdEgd/YcQHvuMvhXKvgolNdXIw5XZ86p45
7rnfCaoXInKo3KVrLeXwn9kVKO4FUufP1+HHU74qBpyx6G7oJq7yB37M0S9eyRDVByadX8u29uDh
5Mrx48EInImJXRpN/UbUUDZtyhDCBVsltbMX1dQKvc+ho1FvXbx8cOrFbEXLH2wN4gwBvNO7Eo+o
dXesrH993xmVztxhU0mxpu+/+HkeWlsdtIc/ZdkfYZs64sWddMw7LR2amDfBzWJfgrwy6y2FNO6z
QU8XddMFjRLIrAUsAgj60dZmNgBVEXI7lZYpSSUEEkAa2vmJ6KsQ26tgPEIk94pC8qTBfKiGYFl8
MJASZX2+N0sWFQ9X/Dngt8LIsl55YN+SyiCS/bEJtd75Wn0359HRyi6A7SN1FVe8SKgZgGMqncNF
2FWDIt+VQD5i2GsnFAM74fI+xj+cf8tc06Q5PeFSftdhNxZe3lm2PRiCqrl7oV4Lh0IewgOtAb+6
IzRrzAg30J+ZtlPdgEOqryU1tNEbTBE+Wege6J5laI9oiJlHI80RT82SAFPw5MqbJx/GSszkPrrm
q3EWnwO2BaIMEJv9mKl7PLOK9xiUblJQWA/FNkqYSVNbsL161nx0iFi0QiWUcUAjfS5++Nfj1W0i
SkacO/GPfv6rhroZUyAx2AftF7HyvVgqoIXUsTbwxyl1ftiP0P4mwDx+OMabgUsFiOww7BKxVN7L
ipTY6sS4PqYeqbQHRFs5l/3ChgTcIWNzQCZWuTM84A5Ocdv7D66TpYvTd5HvL126D33CXXI6e9+J
L8J3XUvU5OouzOmBdB4paO8X1oFFEsimah2a+WRMcWhHMLxQHeAK/WPv5Ja2Vt1p4F2hY/sqEYMA
iCQyc85T0M6oUn+q/ZxSCG4lslJ0reoqbv9QoIwkJpEiq3NLWtNRQb7CUyODfbx6rq4kxAEPmrIJ
Vckv4Xw2VZpYqsl1oriOo5ZulWTQzhc6bjKKrvEEB2PE/w+rGoZ/Y4y/riUUpGFUefy92olvrvIx
e5q20Q0+GjELqYFmVTZOUiwkpXCahtVNylRGHUhunUm/OOJbxdMPxhCGr5Z3sPIi/q/r/qyqgwul
BObsWwfietUJcqkHzKS32SPLnIl4H0yRHdYAFTSHdvf2otyyoJAVMsaU0FjWP5HU6rXNrXLwWclO
KN1Lzh1YMlORykSTSAdg3GbMQ1bFdoVgy5ODmIK+Km7n7kvkGSYVSIrLL/TyrSSQZT90nMjEoghN
dpxd32fLzeAhRBqCh2bQRKG6nB1BWxCOlV0QW05LKwvT3//CAdxnuAfbuk0cu8EWMmtOh1iH9VtF
tXorxR3Xj0GNhM88GnLz5/gF/HId73fGbqeM6rJa2J0jfDsrObAcmqtvmyTvv9hgbo+AXeNBIIux
cHqvYqhX1n2gvTqGfWpWc2y1rybYVQ4tjo89sStmVGAfAtnw9/O3Wn0XFaagyIbQVus6Xo0yVdNm
ywLXWFQ0H96b6kf1groV4agScVd/pBrVwVNS79tasUJhgB1oqSorkLWpJCjzaI4kIy+Zorsr9KSa
GAIqhuVLe3YNpYV53Ud+XqBMpxCUTltazhBfAnE88nCJJ2dSbO5hCkfY0SAC+ObwlVJgaL66pGjC
+uVscG2+p+hnqTIzUEGUoSllr9uWPr3c36iRswGsirhX7HMqc3YHT/S8DguMbzZMvi9iuAGUV4yj
4msMNq+fiJ8ZPBaSJBg7KWbmzlcrJN/ImIX8b/VLh83b+0XCUv3X/1j301Fiq9KTYI/lFP0jMT7a
pURjjvIHzwVZEs6olbtaZmO/cAYAVT7nemuP67fqeLP3r5KZqaM19Iz+v10VVRvk7crUvxeZeM4K
90bgNU2IutE2E3067m5H3Tv7nT1Yb+NpiPMwXAM2Gar4PhWhVHvI4HnEBm1F7sQgd+XKnCvBMydr
W5Jxs/+L954YjLGl1NO6yIVEit2z0Q5B4ag347vGyCloWps4sCHFHiKQb5pikBOuXqzR9iUL43Tz
uR6TMadUQujRLIYC/0vXe9UtyUNYgdOWGZoUtS1B8W7Ky8OZQY7NU4IXZE0IoduOTCIYNoYEDBIe
5alhrcUTf8y5rcYRyCCHivL9FOZvr65tnHahoPVs8bxu4PFpSZ8f96HLm29EFPlCrL76fSuDpmeL
PGkMi2wl1zWB1u7pO//GUeAm1vZ4qYHoXJt51wOlN1NMWvpu/fWlTl3VhqdRCz1izUpw50LcwMI1
j9d1RG1nmgP20tbcYTaKK+ZQgqDqslID+5r6yyaVmeNsOi8ZEpxEejPjF3aC0rXX4ev2KBHs6rE9
1gKyaRlVkO65l7XCmwU7Uzmt4u4zAgdUJyQuTmWMSQGyyMAKM95O3d4tOsCbPqgtAkLAHr3Wyzp9
SmPF6eCRAkH+wPpjDRE/ZtFQzBfNJX69iL17aFRtlps6X491HdyOvIQZXF/k5BhtS0RVWmRTIUSe
YkElO6pY2SjpaUdmP33zmdnBdTRfjsVvEB7fHV4NUxcjLyuIsRY2Kd/TV1YPUP5ry8JqCqLjLvH9
Od4HTfbrQVIPI38MnR5mzvCG/t6FikCMUSGo4oSmjOqan/ea5N7NlL/wQ0B+/5PuFNgD7uXYb1K/
R7jY9BEeE/TykqkjXul4vtPcA2WF+wE/VHB9vp9ID/1+pAQL1pZKlo/KhEEFmiJSO42r3NanKISv
ckdg4v1Vb8is6D7XGOyuhvZ5C25dnYZrOSo17yA1dM9eWY5/K00Dr7310KQrfDwvVC0XQLeTauy6
wVmIHsf7OCskxL8E3SWtSCy/wqrxwFONiCiJ7DKCJvEYoa3NSL7OeTijK8ncs+B2j14Kfny5/iSw
tS1mcO3i3LtRFK1r63Re8urU2aoTV9EsvQ+nfeVqpln7Dyk6W8gadD/tsy+Is6kdASJpIk2gyG6E
kbshbsIHEUo6JV7tjjIBKoaH+liLOYOmFScJRc8tyQyj9iNUtHDUpQKa0lZm1SR6D2vP5bBHXfd2
TP2y/W1deSVaxCBr/CqYi0KZtVac+tba6zENIFUhj+nb3+UW6eY4EQaiFQZOXE93Kn95zj4NCBOk
eZn6KP8ZtXyOKg5t+95rfa6S63QWO0SdSeWZPj3lQFj8aUILnaeUQYrJq0xevTylvRYGsVlNivT6
E3B0VJ4ETg0Thk1eH2Rss/6fBgFsHFgxIuKNXtLXOaUlFSajQzHHa7Ze3PBMeyRWap9LiRDnQutt
GctWUp/Xf55y4DoJe6jImoMfqrmmpNf0FFcz5OOTH5H16c7QD2FuBi7wXgALb/T+e6iRi0zjpdFL
0zeiJtRJnR2DNY95FvnFr1mSpYUGq7dsxYdoiSVrEmIHZB1M2l/C9/GQKC/4Tm0HAhU8sphsnavH
ACIBaOnr+BDO14wiqI/LAyRf63NvetUzqT+jNsosW43iQ8jGvVMZoG+nmMtsm3eNcfKzyHI5LrVr
2+bt7I5lsrG8S6jjcatE7zQkKAY5yoXnubMQWkviETQw2qJiy/kWGlhABw9Hlsrl2//kWHR8EuIn
/7rrbeN2TVfCczZvHNzPQOzrdt60AY15MTOah4o0EXEPaAKdKeGibZrMbY88yqx6b0vbuGlu967O
ECkBLQnbWCV7JIhPSIyU6OeDKyMwxlPhy3MTM/JJyVwQ7TayhTDZ1t+2MTfDD836AXhsOAnUFKEn
Wt7Gf/yMvNDFOPWrnl+iwVkewjpoKaxzu7cZc1KI0Lp2tlyp0P4fpYrxVhpqWjraYpJYSYT+dNXA
KBybo1PqaimMaBRBSOLQj8X2lQuVyJ++Fx8IxLSkxZvTZk84ofZYEG4RdkcLQCKsWdKHZYAbsIAV
WxY24UjJ0lhPNTxNkn8xC2RZJ9/OuiOLoDObsx+F1Bhhq01cVarskd2YLwpe+thdc9YfpgfGFh0W
JCPbpZP6ILuVLjKOK74cgHQqvbOWs3D3uFlK/gcMnzPT5BTB6HabrwK6D+BOV/L829c68iA7wC9D
QWa3j3Gtw7JWT8+mtU0hxED9M0Xic0uamPhXe9HXgVh3yC3xmb152pzthWPU4T6h2kWiHOxl0UIf
Hr6RgRqFcxtEO5/20TGFIDFF5CQY1uO2lXVwA/Vddz7Rm0cECmH3F0S7wCymFTTknBMya2f1ldRH
9HcIwHXQwcJJvYCIFEpcm+0afpMyQ7iNTxzRp8uojDAi/u2Gu6UEUgAwfF7LpLPs1l9CMZsi1AwO
6zdf7EtfB5OClidNixA6RMncem53EJbMJeY/OYx/izl627isCj2nRPxBEfmnO4oA1PgC9soBjrQ9
17NzXtPanBTaod0MQthvgw6eMg5yCD4PTpkV3NlbLqZ4X3+Mcu50H/dl/A7lyAk4Ym0gqHQle+Aa
gLJbHQQDhHjGCWI1tZovl4/odKFieTMACuePSVW4qZZTJqSVmwKDtsSAcUq41W48EiOiboozpUy1
+g2xrcxrrxTlnjXgv25VSxtttjkZaGUTMq8UpLmHwQQCqs2KOWsDgnvxrhsFufv0o7C2ajzrEEua
mKjg3Fg+piw1KWFA7psMwRaDwQ0LHVwt8UMBSlYlrIpH2LKdxmNiH+LhnIhOHDiSwWT4Fi8dmFph
ODwxP7AyR3gj4C9/ZOnqQcejX3pJBZlBqKjwZlcDNJMohA9CjeRlsNhU10Wwr5SElSeKd1Ft8DYY
UcfPWC5loqEidNZz3oF2DXN+bpC5jM/Ld3FYmG+zwQoA7OyS5XkZBEupzSx4/3QcWSB/Wzvu25pc
yXhk9QjFWWLeDlwh1F5yFgJ50BQlSCFjz2Stk5waqxbULWmKwo03Hqflha3g6Dr6HrNvPABqFTCj
4C3HM1gAvd+b3c2yIlpXwfnzepvwnMIf8IsEzGn4xVURRP+KyCurg8pkR5HDs1IoGtg5KiggKye+
Y696TYW5FI/GQJ32wuwt4a//8CeferE6Gomni6XJM9SwXG/rI7v90YZjoEn4zTdO6+0rqmOKRer3
ek1xVtEZaKlyTZ0PFRm7jkU91S3QrILrPqkamCd8pxcZ978ClOIWQwS9pGrBR/hkdGzb0ngEBiBF
G/6qzvfSguv8FvnowWrY/VhhKD3et13XeYdyik3FADSQOHfVPc1udE6kH3zC0mrc8hK4gXVeCjDH
PqGXiGLkzE+/J45yQbNO3vLy885XaK2F5e2f2NhX08Y9rPteLfrCt9iF+fiFrqsN/Kgl52rgtSZo
HHJeneGqGMmMIsBvKpRVJ3okmYmz2q/wmahB+uf8ObcV5lt/5SbAR8MvxUcQUZ9cFNBgcZHh+LpK
7GcrUlq68G4K7k4598PNv1zK3SK8lIX3t4JcZwLpWyQ95KsxbzH5aDPL9QnIdrqCOb8dkWBfd0Jl
cJ4qjlHcHkp7EISzvZ908poLaFD4gjvghizdNFpnxIyNUAIivfEkIU962T4LgfgYhc4h8fuz5Mak
H0+PFoktT1iLA+8xn+ALpR/Z49vHyNCThicOZp61ssPbTKekV3Kvk/H3NdH+rhzsMhrVl9kQDydn
aA85Wrd33uE5i12jx7EVyB1wc1DxYWnVK+qMOnwCet9JaRgVFnV/wxsFqPA5P9zTG3CL6VhPtRCK
/PBchDYNobaV4UtLPnufdEUqDDHnmK4Wk3s562Lh7Id/QF+ZlarSrtJAjpyRbFGsRhTGvMhKgA25
ZLs9INHZjYuu42jtkGYzg+GyZ5sAZQYMN+O90P9xU/yyAMAIa7ymMY/OzU9EnYsdW4nqTXIa3oLd
Kr1sc6m6RsOyTlw6uqLwLA8DDZMug3ONqxyXc9bj3rcLl9Oaf3ipXa9O1Nkpb29GDrcCpkn5Iql5
bLbkromm4HtoUcF1xY+d5lmH22jSAibxorQ5oiec+WLgT4Z312m5c63O5ijcB9H32oWjM+gY7Rov
zJKJ+kZBk7sFvH3N8/Q/Fo1vilqEUpg9NXqFRICwbGywuzcJzdOt2Crts2L1tosuZ9wp2QEHJHnA
uscAuvvgQfKEhr6ClngUrP7/m+7mcYPsJj6TnRk37k+TNe5rYm5g2RFnx6STsddFLmh70TOpJDpN
Qyl8Jsq6uqjlyqeBICSx3ozngUIAT6RUnk6pFMFZbAYcOQQkle0U+0kaMA6U76/3jDHIpLp8OEJA
LUghwJkS4DIikQtAbUKrXXEDSzpK+nJvYBohMxTXO4y35VAJ5sfHceZZ5LsaxB9u7D+HrefmteDK
7ECX5ogmwjQEdfVtOqIwRe8EWVpXZVGVI1rNzwvs7Hv1bmYK8DgVhlMrRsWYYCq5XhFp0ti5IK3b
OfIiLIkFY9xRz1MYMYpSMwZM3FIijB1AvhSi0JUHj+J5fPV8XUw7Rl2lj0ZBRAYUwyJ903buvDAT
5jfP5FmVJ33wSHLEmqtQ2fAPVNj6usxmWt65uXYhQw822xE8t6T5ZbnrqXOXVe9pzEPAJWekgv5x
scu+MKsXtxo1G9bICYX3uR11cGAlrUPS/6PHGSpwBqwaCYt0d1VP/zZJWpVEubMWwrpHSTNpaX4K
3MzA2Sq8cavrhqOEyLwEWr26biNszCXokrmeos5oeyQxINy+WgFHj6ZtbxehDPlSxbUKiYAdbrMR
lO0miJmlcxPjr3wx67lz06XgtY2kTYGQTlD0lEaVncfHrCgz7Vk0/MHVJFZviDQeTmYw4z0q0e6x
IlSOXCTAKlunZJqbkVMLj5Yqsvf2+FI6zwyiUZPVB6tQrDIuuBKpMjt7LhT4nUO352HBINgmcclE
jraATyk67zdkaQUGebvmRdxtkE6zcyuzNaSItmHEt9MeqzQsYWOoGo+zCkexygiztdmfR+84bSZl
a34BQevCscm8S3kuhxiB+7973FX/80BoTFRxKC4Bmpv1TPG7Ubi1FW+UUylZLiOr4i61eWOOd0/7
sjLd36bmyly5C/T4ZXevSP/GQXoDBWzt+3k/0bShgQXdCHEElv4HFVxmdXkZCoMjW+OrxY/YXNZS
LxJUKlOJn0MB/aHNNep0ya1j49SdG5P02d08dPZaziFcQHiRbOwSLxeLcjrRn1k9gPOWgHK1HoVs
bJHbEjLkf8a5rJibRUadWgtxQhvnFbx7V9CoQTSI9UjNEUg6AkkliCvA2geN9jaZWwoqVY5Geh2D
Jsfya127QyQNAMTVkal439PrSLV6o9rL/inGQVL5Na5WxcvgFpamIzNGRiRfga2+pnIbAIjHyBVC
jvZMJvUapx269qX8qRfJ4MGYtcBk8/kB/LtIN/N+j5POCHNXnSSXFSjvIHLlWNhmMOZ60wYbPBCE
BvITAKlx63U9Zf6HgNnpdDLR1gzmONmgdTjkER9NYdog+re9w67Yqi0GSljALseMUpbsHNWEnHwW
ESUGVjxdQhK/E4p0WdW7+HCSirXnXLO4bW7vXCxKgpshpsfIRoXiPBr8PbH3yzPXpZrRs7pC9Kqb
CMEGxOFgABegzkuizuMa8jZHRC3TDQQs939QkqZC7zMlnvKanwy+B6DdVjB6jIt32NC6iNDfKaUl
9ZCj7EVyDyVb6emjXky5X7GUvKqpHbKi9N5aNaU+tDwLMwCy6qonfCtId5o+huGngXZhT0DT6L3O
eMmRmxPezl7bwSTojmf0lQAW4iXri+Rg4my/zpN/JXSYAcidTam7HsEZjnx0+VnB3E5vedeYEENO
ZkUHcyIzu/rHev8Dg2o1kw0LXs8iq5I0dh+KU0SkOWCT9HYp7sYxkq4mzptVriM4rCOruPghspWh
2PW50Jp/TCEeVVRYmiWT90aszSUZGF75Llnl0l3xZwUauL8w2NrRgfFH1dM/I8h5DW/e7eVWJjBt
TvxhZiWdMgcWmax13ihcowOi3og4N6vHupxuYoDWaRM+aJJ+oEeN43MXJLJzyNrpP8yyWoM+29NF
n46KVogcYPs+RqVipnNUi6anp1glvQ81aDMxN5t/P1oDxyZ+FGvVE7Pw3xvT8RE0s2A6vd8f9JF+
p8CgWNiF3zCrMgvTe1S/sLJ7N6NrPmcYgcCuDVmfQ1+xp8JB0bIEfnMBC19a4ZLfeUX8nHbGxZ/g
qDqRTbSCtHYjlbRFctvxoqClgZRscwymAG80ni5W3SEWGmA7cfG5UX6SVsHzi9vsGUgOpe5YgRUh
EscSymRWwadGiivEX19ZZvYEZrCOJCGh+WR0uzuY6Bh2QhUiw94LA/w8b1XkTO9oFILQ1OaZr0ex
OoTGKK1qqo59XUZWGn4w0fSUhWcyl7ZZZkfBtbQnyY7WuPENZ1D9X7TnjGBQUpayQWlixe/Dmr1B
PMC/qH+qhtfrdcTE9A0jkxzwfx77txHTOrQ3/OCmPOyHee9CXyWHm41dNM5rdnlWkmvgKB+G6gIY
9YRzeSyEI2Qet2AxyMO7xwgEQiNYwMtoh42C1oOfTndnk5Xr5EHBVpgZxG9sSzzwiNmNhSVzBC9L
xCBfypypR9lQWaLYfMfG4tgB0EX2q8GBDwSYWt3HOGv/RPItID5cPP6anK2M12vzCiZGv/gUlKJP
sZTUOPWO+wS4wHbZ0gPnZq2Ltweu9OY6eKz9MSsPXyaMNvH/aPH6AqA9Yc4JiHhIkAS4mcklE/hq
36FpCwLO6BPwcNUR1laFUss1w8Zv/5Hn8RHa5SoAUruH+kwSMZFT1o+jjq63mnvX+wQcvSdwwkn6
X4RhpNvwwBcTgbME0ZRCOWRl9WAMiC6WtTMfAIDvQlWxKaKnKsZg+0OXglEMe3epHVAoawIqJwNE
QiBzWdzdubkvBR814pRanutHDH3WUKvhSb9sPR9tYZ8fTJ4TmPJ2fJ34IubCrEWBPDUA670WzIwE
YqvAbD+qpTTytp250NLGwHpXz+SxPo+1ITRCYpAPHVhmXcjQ4R2mPxgkVfxGLg1eRiyNNMUNzSuG
oxSMODYeNBLTlN21qz3x2lf//VCWUgR8v72FmIyOcQexIFcJr8P2YHkTNTjcq96V5BkQ0SYd7C83
PXLSz0ylF3ySpDFRgs7SwAYGYW/8pvvGTUrQt3cfp/926JH9QXS1Z7GQ0MxpTCCaR93ltHRSLfX/
+u1oNvcRgyKqY8/U6M9VV7PzENbflZui0gQUqnH32emXhYPkhC9GIe9iBWQjgyH7Z8oNL9Oskz4B
+16X0qGwbyNtycKml2T86r87gsjYmlM/zrWC9fEGnKbr15xzJave8clb24d7YwRW5nbt9hK3HFU6
RJ0IgjM2urQD/lEspq0rhylplZeaObR8i3CLwe7teF0ZR7N7xeQSxsqMDCUAgWxEAUzH8olwS5H0
3nKd341oNmt6NpTT65Gy6Oy6kW0hazL6ajhszPY1g2hxbAnflfGoT1Ss+/22dh4u3Vf1uqecMOaO
5faBsijUZW5I8S47HGRMUIffaQgDaOUBbcNliWKBuyv8f2LQecsJMi4RJHc51Qo/zZEcNIUn5nEt
2lD7wtDRz14GudClDPYJsF75iKQpyJJ1zOukqR4rKfzOflAaNenyDiMUXBuvQh+PxgEX9ua/UQjd
rVI7atYdrCJ/heJmS83E3YWireNcZJFWxQNNpqwcRFdsIY20YNQkjgPiHpsuUeHL/PW8LSKPBs6t
Z/5SaWAUYsIopf3bPw0LbXUXu5esa0WTv7dJayC+ziHTLJ72z28HNsRHP80c8dBnxJZ4NtSPg4V6
GjH1GxGCLqEBxrn+zNMInGd7K03mDOMv+k7l8RtL3wjnm/C37BBukEEEHpJWPkjJqC9vjtiHpjRD
YGbCz22C06Y5S6pqrdnsP6Uf+UxZ8M/7mQ8BGOJj6N5X9HBcRcpQCMzV5jgj8Pm/dZLQpZU4qIcQ
F7meQJPKigeTyD9TrNqS2p3HNgtVsAOwIsWnIzyLkQPPaGKL3+xlxTQV5oV9w29i1dkdwcqJkhCE
KqKb9zCMUfH9fIRvI9ymu5M+rMtNkLlKUnLja7E8rMheZ3OoJviFiv+6DPc2IQuc44pUs0u2PiAQ
qswfbIvBA/Mh/y7YObqzQSQ10DjEyA9KwUszHkuawSL/222Mwhls4zHZARuw9FAkwiY6hiBLrmwq
vB0XPuPSjFcYAggj79vw7Gc5wsXtfv5n/qU4eqKF78fqqvh+G9JxjT7YHO4HXDVPTWnn9vnV974J
td9e+5fn7WScgvYok8EXa7IXGvs3Wb4AyH7KveESMN7LtUfXlKAj96VHX7st0GTJfPTZJGW+5doT
UssqOdyKe5HKD6KiLGimSgZGkBJaXDEqxZyDVCGQxeqIVDIDKKUcmfN7GQcURpWj2AckWJPyfFIf
GLyHYDZiZfffg58bvNPFgiYR+vI6/B93dXhzamDKt3kX08QJAdLMsujIXFgp4IWtBOVd28/GCFc5
9Cq8RJhhZYWxfBv2SbXsDQckdlRCYkB2iw6dTEJyTlpnR2dsWSMjhsWD60F68rfwzP6FFiU0bx8I
euvX2tbc63WX/VlPn8KdNMBxvnr7VdO1XXHcVGSyM19QlrCXHPUSgbYFEj7IPAdUv7R/AZo/C/Sc
hvDWx5ZUr9HiuD2R81PmtDIlarDDchOG2rD6S0I34zRUuTkVaN8D4NsFnvVNR3cUoWylfEAckk8/
xI+1UJi4AlvKESOyDLtfAfu+uC8xOU1azWG7UqTVShhW6QYHBwiq18TL08yFcpHCWnPrhbzRA/8V
ZFN5x3MG+ksAGX1jzw1B1ktNCLX0K4Mz987M2rH17PPk9Ra/ZKduwkUcr2e7U8LXdurpmUN8kjBM
WD1ggWKF3cAEurqFu9KFCHiHOzvL0Lq+HGCPqtxRN9XsItExWF3z/0Zj1OqTM8fxdXB6SzART3mq
KqVbmBQgICPNjWjXl0E7Lcb9PcgwKYTHNEWhIdvsFu4MzahXGDeZxwChfTcvrFgs0bmCgS4hkgyQ
TtDt4L24EzMqJpBazV9XdTlewsg4rV7ybPkQLfq+dfiunwKNVxhlMpMwI/e8wr17tctcwvS1mfdf
FWu37FzzNVidZKyRGasrb/hmadhOMF1TogDzetTdM1rHOlZQwdwh4Nn/IusYzvsf3C7qh9Hgl4os
rvmV+6qXDd0lm9TkYj6PKXtgFsNaITUpZgqwC9O13OflEuP7+qEeZlpDBda9I3fo1Yjq8GLRXLvr
LUmOnFtLC3+bBFcvSPIU7/LX4YtZXRU9rjuK1rBJBF6cDPYPgVPM4b5BxI4GxDeswdUlppz7GGTs
vgDxdQxxX1rvzqLCoywfRUAHbf3EIC7LfuLUQNXGNXzHZfZx6GON1eJRcv8gcTaSfMWhuMIvmH8u
c/NRZDokZW2kqr2YT9iM/YSyxsnih0pZ4Ogn48+CcLcFfNIHKkuu4fkoamaAoZWqTHWTQStgLsYD
V2DkjnobprX5Fq2ij612/M/W3+gt9fFjxbcHQ1lN/DV4Yppmw4gEqMf4rLU+7wRFxh4QgTxO6Jts
GjIvu5cIEAaFASOP3AMkRsGNu+qR3rQzQ6I0g8gr3iWZuTKwU/MdErgMuK1v+yY8sOEbjPeqxxA7
131QkgNPK/wGgOFTaUcIfO8jVt+HsF6REQwjjNF/W8/uziAAsWCH6qKUtrcIyhwyCV2QxYEDAYzw
x232mRoFqGrFNaXM5IVO3EXbGngwJuJ9cc4y08vq0dSgbUCxk0ItZUJTdbWn1e7hSGkf9zs4IJHx
UmjXTpEKMrZuNkQo7QWV3U3ykHohxp/wl1h+SFkQT3Yo14kzT1QZZVy2eBJGDB3oVIpJ9p4FKxfm
VHS9QjqESDOSqPHqcJ6HahwkgtTeHsHD0LOufhRzTDJT1lWuegknf65s/JJ2CmCe/QQYfkRYqGTo
2k2uAlKEZvgE+nSzbh25rdrhhc0Ds/ezoHqzsGbiL8+EUQJUA6BSBMfqizikuuHnyXaOc47nuW+s
m9fCNyzCBX/2glJJIhOYnaPuPXdvraWr6NYH8UazvyzSz6QFQml0Hz/E+43ASALq5Ppga/OHexP+
887yappsMr2R8yNULVpbfsjWVq4TVzbOVEj1BuivH15MV06SN73EZXJHSr3JQNQiEvKJA0xGJmCW
C5Dr30ciU/lX0AnERSmQxeM3oyC+zzHGhvOUeUnI1eUsgh91p+f0Kh8osKadEOX/xrO0T/9PZ1UG
ZrYuYxb73wZPwMXxNgMJ37c3PnJ46Kvluhz9dzdSuo15tDJlUVR6amOSSi73ATe8Z+9VaxI3xyN3
2I+Lgq9GrlhF8zB7+azWcZGELgSFENx+UC3YcQteVI8uYiL9qNeDZNtilOG8vpi12q3wlQ2UQvP2
rpEtY0Q2SwQEbQWzbQ1wZ4NoB9FjuAKTRXpHX4aRdtxWk1qDlFnlswCvtLSbg4pbk3UU89+GpJ1D
F4AJCfbvfyo72rE2wwMsRn/wYmq3q8xeOx18PiAkJv04QR+bxUG85thKkfmDmv4GCMvM26R8BljB
yM+B+SyZ8OI7y55/J70QHtbIlno7AK+1puAKxCwgCpcscyRTx6X+yNlWxs7D3IBCipJ7FZk29oe5
ahG2glahWJhgX1pUVjz7FHce1smwtVY0R9dceOIgpUBwrVhnRaE0fa84GX7dBHg17mHfzemZ7hWq
5jcwcx/kv49tDGeu5OMi8QVYRuD1IsF8tHLPrvGAXiGttfSHT749TxvEjx14VAyGp/Gmni5ZuO94
y6thgXz6aUwnsdqayOCjf+1hc+pCPtU2AYX32oGwvzJMIBwOFqLpc1JR818Usaam4Pa1hFaPaOfj
riQMA/9Nq8+2TVyZ5Ft/XLgq6443zX2MKpNu9JKTT6Ui2Fw15WrQzcFYRN1tV5s/yFLg4V/dlFmW
5tBAs9x6mdX2d+s5VGySLEJLiv/JNY+5Sefnw5bGvswnthgiiAgoQvuuCu24RUMCxhKHPgiYCkUm
9bSmX+Ilw0Mp1Um8q9XVCfjSMYbCjSNIbesZrET58aGCObRATF88yMv/4MjiHy+N+O19L9KBpPgS
yzMvvol8AL3Hin0SHPG2gSc2Kfg8xqY2ICtnXgsdi+H7NBhFSFfqXy4Tt7/oNVwfBDrpSqY/qT/h
MeFzvBwo5yXBPaa/shBE01ylYjZZEXvCmpfQ4b2tLy9S9ZSoFsAbU4vMVwJYxCTfXixuWD915c/Y
qfK9XWrWZyqEDgorVIP3n2W54KrK5IvDRIAmfvC0XOfA5QvrswxVgoKnCE5j7MGNs853SEp/Hg+u
7u/HSHkN4KXy0+5CKO16jnxof+ooxBOC1gFf+ke/rNFzfLrVjFU5DNkMMhY7b6Z/tfgDLeTAKZtZ
AY3YM1dVTsZlfrNEMwo9dSkGNgzaxwDjDi6TbE4uJ2OUBe/xhcQP5/CA/C2YpT38euRprtfllbyY
kXvOtHuZAqGAVCUisyFIm77acetD45RjORiwe159gxDjwJsxcv45/pjydKv6BmjKj2t81vhjMdFR
72FHJ/XrTvH5PO6FQ60ENJtqRnqb1oRwCD1gn0tSMXLJ/8FWyqOBzb5G1AML29W4w7lZBXp3bQxB
BpoOs+fuR7r4SQjIcHMVedOcocENqyevGFsD21Gy3FY0FKWOqchfeVCKTYMLjb41i9ktp9w8G7Ps
1txUwpqkc2Qkqo++/sr8iAKTAPMhcoe5JwS+FWo4/jhlgpZ0Vt+ko5rLN/Kn9/jVWbcaIkACfb7s
231y4crFmCS+xzaFj6Lzbk+scPp3STwNfT2OsTMgIY7TbOGf0AzsbYfYO1UPx6QfWiqMMylFjPCR
cvw0FH5a9jPoNo+12JHA7gz2OUL87Emj+vpxGZNvZtj8Sqfp+m06jeT0whG7X1zgC3WpHvIMIUCR
P11BxhvquhgRHFTH4lg0BN5GrDsHUEf4e8XYyzJ5o0IOj2hxCzN9Pb8LBES4a3N7ELHpuMnA5Yk0
EAibtFpeZ94DxOTG04u1UAnNDvGx8m+0sw2ycIf+lfQfKM49tYhjVDxISjuAEqbLxDksXcLe1Uyu
YYRi7Y+fSHBF6IjjrVqHG24K9ULJu+36OlHmjZrsY2ecmCQkjf5hpemsEUpvGWXCnT1012XtwEMa
krAbRCTzZBE7osG75nehtolSoIuUlIQ6QlKbl4vxBM4VOufg+6mxPagDhE1bpWviCo0KO9DCiygx
zncNUamkeIGpzZNix+NnCmZ8OSBLNeBaZZwgbPGYFS/FYkXegJbUz10lGQILUXq++J/k1Q4smdFx
P+6kU4QLz7YN49k+REfSGU3f8qCSIqX02oxT2CCVsaFEgAddW9wqbRzQcr8awzzYjAMcufBAsmZa
gZw9a8OzNRD42gkrlteUCHDAIhaE2T1pcZsXW509sntA1TQhlyDScv+zVXHw2l92WQgsfrGRhpHP
DqJrO50Zy5y13U6pnOBhZjPfgsRLxS5Lz1E1S68VkH2wLi1oJASR7VMTbL28SnXiQw7xf42AzuN8
HJi/IpOpV4cD01NxUWcsWaUTbIYcchFn9aJCqPGAmieApTSKS2Yz522JW5i5hX+3Tk0ejjhyor0U
Zji9jQQ+wEvUMKRhf6GDhETTh6ctt4pugVvbirvsNYgoqNPJvb55z7hsybi3NWMsO61RYyis9/Qw
tw0MipBzgA3C5u/MgnBHadwBkFSH1XT/vih6enNTig1u45MIfxDJYnY/2wRxIr5FR7Ezz3jfOaGu
ubwFyXFuWpiWQjBspkCi1uuajuCXp64ZYCgukVh5r+k5MULC7iw4tWsW6vdWIPS8IRo/pN4HikWZ
BALlDg/TtpB9N2K2ByEIyElmmYF2OQndIvoq9veghfmLijBh+jnYPgvz2bHFvUjkUsXW/RKuT6bQ
w12YaxoHlhhqJv8AIMMUT3btTJOb2nRTImrA2dSJtZ5SPgCnomKF8JjQmGpxpchRoFBon8UXmb6k
2zSy3Cb03d9Ra38A5Kwtr1cZz5aoV4Zx4QZQtGZSTqMLPxDfYv5X1N2E9yDhtFFHBYCUQ11nSyOB
Y0P/5ijgEcP3vuddAVV4uz/TT/AMJTCjCophpE/bjWCrgvLcogPtw7OoFimwFIJAJDgN0Vn1fLVa
UMY865+x1AI17uAaFD/P9AGFUhnuWl4okbc4kacCrDQbr3zQFTxn7RiQq0FYzaQPSeDkXHBgqH9a
jcOCEAyJqoYgZL+A0y28i73GcyTgFAoriXp7NszJIujnBL6fNxjQcrM3KWZSRsX+whu+tkGxqG29
C4ktyi/AvZrcfyLC+0GjC5+Q+Rh3UGQXLS5aMadj8M2NzPEsl6XjEePg03q6AnJe4X8jqlPzCO91
eMhzQpC40o5GLjJ8EMrEmfNr0+kYxRPxcqi7qInFtILvZbBUaPTRm464/MkBEzl41bSyowhwM1wL
N+c9w/LT81x6QJgfyFtmglC0VrC5+9zX1WIAieMO1LXtsQOOLbSZg80uyDAzoLMc5LGF2+mVWzDi
+GIgPtvtJPeRsShvapj/6+G6jPbvQccEsTlLDA+M2nOjmmhSpUlcRXGq7uBZqetUIXnMBLcijHV3
Wg2ijksVuiiom6w/5jdkNABBwPr4lvfq4I5RxY27g/BX066CkbOXdhRUm6mGaBVfDVgAlfpQ92yx
o7BnRa9zYpCVFw20OmJbblopgfmuX9bK0O3NupS03TOtflUTFF8qb5Hr4kOHdoXtf40fbUtFEjXu
zTRDg6wkq7TZryErSAVqhewqxQj5wcSyOABnIg3PFVDCGO6urniCwEnWZl/7VrCB1K+AQqYh0zbs
G75Dl91JLfMCOlxvSDFAeWosfUsid5I1+MvAATFJTxSP5OYm9Rv6ygz0Mo/JbnkwpuSIrugsMI/x
p74GlwxCE+0OejupIJDipv3UycM2joZNR5tIRsWIzRaSDBoPXK8ym9eS9B5TuJxvwBInAunVlyfm
BpFc++WRVKBsseFMNTJybL72e+3wLCzJ2/t04SYX0QSVJwysS0s6DCaUQ5rGOzB8j3AZcCg4zg2w
vGdgkZ/t/dMVPdsPg0T1Ogb92tBssy3S7AfcJHp0TVWQYBSfjpSWIu7d2U6K1/wYAeLeDvJzUsA8
DWOe5kjvIrS9Nn5wZP69Y2JU7ZysLFIshhpPFvsE3Mw5MawDUJnlfF6cXSJY72Ty8IgnyB2krmsU
qDE+lXR6sRfJZ3FGfjAyVjDKMEXiuYEM9ZOTEiDqFq3iWINlaYj7UuPs7sV/r+l1YnVTANLatrhC
0S/937d8xtd10RmxpDMTjb0WE0UCxlIB6SQkqzSIj5SHowydKgPEqO7J+WupsyPl/SA0HIqToN5Y
Y7W8xO0/7SM5Y6ZOPBYeT93xzkDuTwpPXgdL5xpl7BgeZBc9rD0QxU0qGgjiszB7YywpoE05Eapl
6c4rxlzvpojXDdWL68a1YJj60KWswby7XfuyrT7upzR8DTvhY2udCcDS9xC2E5bYDWiosprwiTSk
UHwap2QAAUmasAl3pvv+FOajycthWOtWJQkwjnNuj3KI4Anyr9191eCBMxm+8Pc0VoLVz3X2xKxr
9ucuPTD4CsMBKP23luxZjRjCaGdCr1rG6aNZVLoQc8Y1IuPH5R4z0TjIas7r5LUayP5h+kBAfSYS
to2q9V+fEdtH5YmF7atPsgeX/jMRzPQ+yCHUcPTSidgidt4vh1GOJS7oIZctDwpcBDS7vSIB8SRo
Fyg051yQJQ6kz3E4Ct5s0nkS5JZgOB0JgQz15qKvnDiAwRTKBHFI/wdHyTVowdoXN25jIY+c3eVA
cHfEuiPXkupILEhIOErPpmHF5XMWqBlPX7tIt3D/XOJbPCroThkWGcywNadWg4bUFIQyII0ikGFf
dOq/W3gUNk868/QppnJ7T6XA/KX67qLTbjC4YHeOF7rrvIcw7QytNliIQf+jWmRTrMvZL/fzBo/a
zlo2UI0oKMS7o3WLRtsaf/NBebUBP3hnKTwL3OAI3h+dAUG/rb+OicGKpUXTA5fqmTHWG82W8YGv
M7wIkBIjoptUINI0taP2vxwcKb7SZcJYed+kEqx5L+f+SpfOomzmxQInTynubWjMSzC9Cb2MPuAY
ooI2sBjVogbp/tZwKNRwRKdhb8JVgpKDnKvBY4tWUIyiIoNvF9NhfiUYFRzk1x0aA3gPsOvIN6e7
8T5dWrBPRvMLJZjqy6CFK8uN3m9pysBxkgslD9EZ8n9Qi2xMtWC90wEvahOIJ2++oPXNUYGzpi6g
uS8nAUMwaAVDutvtKMs0yE23uyLIlai3iCbHFi3dEpa7iU+G1nT0alCxO/wf38LqKeFKt3cH4f0f
0OShxXcSw9I5U5tH2XpMc/5xwdK4Snj+IQ/Kl1kWO9DDotuvz3aVDr0ziQlAuMcldOiAkTjZ1xry
4UhB7xcU5EByw47CnF3BvNYCPpkUBQH9O8dZjnZ3Qx6EZevtmMN1aoIaUcsp8dI8vANumL7ATVXU
gqDTnfSKMZpO++57u5uMWNCb7igA0d5cFzalO4bJxNPiegwwMlnfbdggAWJdaHkx/k9NcRDaAvOA
QZk4fJPqd0GvSSgr8EegqPymg37wF3wE+gD1Syf8i3yeeS/45XLTmH0yuz+o3PGW+OPis6XQV0Sb
c54wD+8Mq6C/e3aZqwSW73CSG2HYMMp7nzIqSjvvEsV3m4kno0ObOTWqLCA2TRJ7ZrpSvFJ1f4rt
bv7uBWZRRtG3Fe4W2gPxWHf42+LcON5XFtBAH3gq7nasO1YkqzVy4IMpWAlkP24N7F2P5pVyZOKi
knR1Nkg8tATRvOFWpRLr0RTiSR3qiHZk1dx2Lu0c6F+0eYwZ+jgIOxj3d6aaVCRsjs5tDSqXw+yE
JJ6tV56KmKwfqytH3pGCCt2tw7V8YB245kdMTVe46Dn4bcBHgk5T1VP7UEKPFW/E+yJSVEriQ7Dh
tCte7ctqgmdAKiXxoeKdok1rSWT5zIfyParBYuQdT37cEMZI7QJf6V7JTZtiLKfgA/WEMbxiBH39
DW6ESK9D/dVxmmq/MiphJQ7EPc9q5LhOJH56X5Pu7TAjYvbSTJy0VefGy6S3fkeSkHD3lSRfOxEp
vYYUS3y7zTVP8rmGGjvfv0msxxTzEk+BF0s4aztTRTgqqkf2h5HmiS4HPDDoLyBxGZi1nRJxsc2/
9D6ow3YLv4J4ll2GTG4Pr/vpFfy+x2LKxN2bFKQ2I/QsmmdJ33cFjblaBUNJkz09e69j6xKEKyKv
SewjwuD36srz/DA2M01f+JghJ8hrY/LhENFlzF32uXOjmakhxWgYAmXO03SGvVK2zBAkn8jCre1E
U+MQ/fzLSzYbvpIP5zzngHtOctYnGPtP5xL5QWS2qniJYW9AviuqTShVAautaKa4p9vzPFLQMyHg
KhvRZbc+xsJhc1ok4lm4hxfNFD+/uWMVlmWxC0EaOZhengWI7x2+9ho3kHP+9ID8zyIXu4teJnc8
vsvA/ax9mb2YyX/W9BW43Drmz829BABOtHulxqLmckVyOZriaJj8QC1PQJcV/RafaIO2tYfa6TjS
QIJ0AK3M4iDZBLKpmQXtrDGSV6RYuysVq6si8hFGWZBM0e3ramzXwIHpn9GnhBEyW7xCQGR8dc5V
zXcm65Sprw4/GgpGsze91m8uu+XS9DBcX3n4iQ8DrOIW6Mdx1j/u5LBmDxmjld9D16wKRwRobpCm
zv6yxY8oLoykF9okfDIbXLtOEsMGVOjrudck1eT1I7aiLIwTg85NWeP7tj1MYNOzBigM+GX0dTtC
3FPPj5X41/SMazBJhAgMwHhDmvdh5e2Ie65XpJWGw+y51C9l67xm4wv21bFCAJrtuUKvO2SQlNyQ
hfoevCvQjGby4COL7OE4bLzpgnBBPlujmsPY/oQFR8lDSBuPSaWj+drLIa+Q4wHpzmL9i9MWjwpq
UJ4Lw5dDCwEJhlvTXIJJH/H8E/ptBcsS0DC66BvxQdtfh/OJwRCXLUqKgMhTe6WH5UzW/JCez3SH
HOgItGPfuhsLmS53r9jBn2CuOyHEANFCAGvt86QIx/Yp6loZFgWFRrJzLYCDCnfS7BFjKwkjSARW
C9KQmHf30d7kc4kOBRIpe37GaQVQ3ICdpSSQz7aPo0Rctngx9e7sjCCm9kDzzXA0EGt86lD7dxUS
HnVzC46OuBx1INLlcnKSxZHBtl05YoCwsVhiwLFI4Ol8gzzX3ybXWMNC9gWjSIAjDJrfen3NEiBW
qqMUSaBYBqIHY/3i/fBvDhzmasO7pB1Y9E+gW7ORWxoza8oEgBR0xFJmjFVEOw7nLzNVAzTHx/Y8
iLU6UiuvK1DyU57jMffofU7gJkhntVLJ5EoHYlQky06Se6dYvQa1ln4Y+Nlp0Typ+yRShy1rgAnF
2qo2pXbAxwZqyesecV84F1tuDosXCa9zLu4a7ZHk0jFpFwGfA9ox+GYpEbD242Cs2GjOwDWnx9XX
tP6gpQOu5/DUyT1p4FztU+5eF6uwKfLMEwu9XIes8Ek1rlSVDdTorAaaAyjIwdSyF9OZ4ZGGKctr
/uSIREXoOzgnBH5R+r3kwgw5/1emdZ+PNOSJzRX2SEyKzkjwsEm3Tg1tXJYooNgBIiKtveVBzUno
9Y6jLMycXXJ3JxzxDzlYaW9rl04eDKSjhgzqWpMxVS582SJfmiHnLvGEsabXSW6GRLTNkuXcnFqn
NUlYRcIMMk17HCkJh0A12vhJkpDCB/W7wtdoEm45WyHZ5MtFsKL/Rlx/umZFk71iPWJdpgwmD331
irHN+iC+jV0chdQXprUxg7b5sPHo6yuz5YNQzr9/aCwtwjfpekWBho+G4dtv8PrbHSb7ccBvT/vz
KWHdBM5Wyux+u0kE8irWh4dyqxJIxWr91bkftXrrgN5chuvaLVtUSncU5vwAi9c1/z7CeM3enf2+
ztA9hfQRYPxXxjsfJo9VxiMipyG9XADdrDGk1Z5Nudf5Yh/bKBigD05VijmCg9CQRyake48dOpHP
Edlz1SM3ZlGiSsCdKnQr5/kJhwaafuZllQmkoHtytiSeMDrDo1OgeFSpsOeUaAvVkowntaOhEWVh
Xvt2UKdYcDVdygnQ0+ALVU6NMpACoIvI+UixOhQJBUaE2HSYVXXC4MwcCFrl+A2Yo35sl3Npc3Z7
R+ZWIWU7RnkyPVLrtizmx41MzCrohF98uC6uAS3Wunm30jPpLc7dVK6rxJnLH7aCONvepg44QBSN
aVKCjEd9De0lXdgWnRqAGNfTBt6WXT3ECCU4hL4UjpsCpNV9lIL0gSL9dSy+ZqPFu8dtOwBm4lBZ
q8EOdx0dSiZKH75xYrZ2M++UtiCFHko2407yvJYSH0lUq1f5YM06TTFj8i88QwhhwAaEG4MlaT3e
ufBmG7/hyt0/bocStAay/7zJQpxs982PF1o4z9w7QtPVkZmm1n/m/QxXXtL+0eFW3kXxsc3v+bqq
Ddsh/22ODgIOdcEi05CHxz+98WCJx7L2gyrKqFqAu3uZgNwV8BKNTbyA8UoWwnowHjbPPDyV8WH9
42TKNn2NtDGhvPzAe2grlL4/1sqTASe1rQL8yupRbTiWTE0DxtTDf1cnc7J/AeJonYgDhFU6cwyZ
GmOpmWGA3prieVrCxJuUf+pfRmJKAD43p16KYAyTiUn2WNL1cfUMtRpfH5WZ6x8fC7V2Wa2f0i7N
k0DX5OrKAQ+iceJpRg6d+niqfcrOygfw35mpLu4PSKfT912P5CptJ4kP7QkQTD/7EcT9Vt4I7Dd3
CsNQL6Cla1Donl8V+A3JTEXtqwo9tCtX89aMU+Jsd5XLkO1QVDyRirLAsqZvqb+FXf6wlxH5xJB1
T4fs8A6dnaH4qrrsXJAxRC678196r+FZcNil6WE5HvA6mIvua/ua61OkOlf8O8FSo16wMf998eUM
YebArTTqkCi074Z4nhQYUxOaGPw3z/cVnrPcDKvH0xLSnHIOMg8VYvb2kJ/gFwauGDWCPhOlVw9M
SBiBEMYttNiStHpOPAwbwcfuAf/W3q4uWGk9EoYNpKekbSKlhmr6sxVJFGxcCzh4XX4z9wiV0xhW
JWJzLXUbbDnX9W0AzYhTRLRZslUJ/F+5MCrBH7uLWg6Jvi7eQhFqj+C/UbssPpwxXzg8HKrYU1QC
MsgsYoxd7dsHN01L/Yq+gO9t+ftcsuHG7g97bfrNdwqMghTh1MSdgkHSdK/PaL5xKcItfdL6Zx/s
gAl/RYQHYF45o8Uf/5waugBFi4dUjxCO/p/gPH3c2dCbqNlGvWG/cTink+Su5O3fGW395C2jeEWc
Bpr6GNOTSvwBf8DfQ8iDAkbTHbAa+hO/czQfgBHI3j5XEBE9ZtUaRIcaXDEbQoLAPxR1ld/GveEq
PEjDUFrQ2iujn+rsvxAdahUqgR5NkcSdgd61aUQ/C0wVVm2gbBxACOyhWWJNJExWr7/mpg0Ed2cl
RpEYSPdsIyzDOjeB0oc2cE3ADFB7vvFjnlBikySf7GtipiVb326cGvCspzRw3Kcbb45GL9sU1Or6
Dx7on9HOmtIam9IWfAW6WKCZOLXo6oWu/VuXaeYh8uibobcq3aCMW3tBHGs7PeVS+GQtRl2kRMbx
TbAPwj96vXZi9+8uPCPSwUz/VCMfdKV/XYgpOcexsTa8rDh6i2yQjC8mrwmBoAcneEFPx0fcytPw
G8+QnTpaDllreg5xm6vBy+lMItFNQ5qSSJ9Vf6SfGsKWSZadWtcg7CwQ1F+LgPWiCawvZ8uxVpSB
nkSsLkw3h94qCOtqnIZlImC6Kw/o7On1VvlAtL6nfD847saE1xYi3c8Xz4SbbeUqUlubF5Hy7gPe
LGTwAbifFLARR+GFSaUZQ+DbI5fSjtyFvI3KVDKZt1gkjd1WujZ1yHACE9/OFVzmiORgg4dRQeJm
FR9RVIduvh3Ld/ICAiytw8ra5/x6PZBA0YyBA8ZtzJx7FThP8nG38i5b2b9z4gIee+DN83e6/eWi
bed3m8lNqF96ihopa3KfABrdwATxOPko5VXADPY6VkNqcOytcMPbAmkD8/nbj6XopgXgxFiVkDyk
sTf+pDpuj27RJpEeaagwWUvqkOf60BXgxxJiGLE7G3Hbtc0TWvYCwtJaZgXkhb9VKYj48/m2KP9/
kIDswgFJRm8fvOdazxawQvvMCpOPAUTxWPiHe0zb2HVrg/kwcCwdMIifmjVvYj6oLBohv8TokfjD
MKSGTEXMF7U9ad6564RgALR9+0HncAPxtdMKewqV3XM1GYR9KZFzcJwHL9+PRFkxUVl83XeRcvvl
xdwsdj6HddtDBiHeeKW1X3wz88EQkhF5N30h9pAoqXHDibHSjIQbHXjN1Hm0a32castllG0ZYxBQ
hmKyIGJEdojWMusDOsSYpHbAntqfeMEF0Z5gBROIFvd1F/AWg3HPTsxwfhfOpI1nrU81q/WMXGYo
DWnST5ELxk6V9uOzVUHWjCh3uX8xl333cU58OUZltL4Tb2ZgPlHQK+DVfw4WrLif31afst8Vfa69
lGXc5WXL8lm+LnBCIxUqV8Ye9jCsZxP/t39wWCaAg26gTu/Vej/6JJVBYeWWhBHiAp1Jo+oafmHN
SFOK0S4Tzs4jSUnl5FEl7Aks8zHdbA2UEH+lm9vKun/OxwS1yJu0h6cIIjYQqfvW69MlEBLfgtI+
kqgZkcjghACX+e2rL42zPDqsZKJ7OiCsa4k5ExT0EIbHfTLHisEDrVcM0SSwwmlLttKgxHRsIWQy
Qiux9ehoSeVaPFSrIzOxX/Qp2mpLjR+Eg6AGXWnJZOp6md3xhEFJ89/bk/TGb7+0cSv2oKImUCLy
UO7QMrkESlHc1UmPP/wWLe03Rb8tpAP4cjWXg4VutLHinS9Lql+tk6NLyXo7+EsL4jTcaceCXGco
kPHVPjVL2NU3qrjKJBfwPRU9ylnW5JbrLqksjoxOcgkYE4ROreC+1jnk8iE2jC+kLsECg/essvRd
ux4pqJrJePGl362qxKS343Q0YlJsoQbrsrTiqlXEjOzWmjYxbbXf3Mlfy7PqWbEfOgdeLQBz/7yf
B4a2v2gOF3xJM2xYqdB2swnEMmml9Y6XLS3uSn8fUdygBplsUmU7uOsMTBb23n7MjaGkEcJG2YAq
Q+AgtCEJlXmDH+kcLP5RLhAu2n6nyBWxIfWtC1tBYnGAu0AQAcBveQ8kzcUmtrj11FLJ6P+36s63
+OW2cDOTUFPO82MfyZnamR37S1V0V9OdfJ+r1UFZB/2SfHSfaekk/d8Q9evAjK7JcHyz6vHY2cNQ
gcNtOhp7yLJeqC9ZKqnefnNd1QvluUwhB3cvJs0GUJk8+uT2e0k665Heqi2wp7GX4hN5Lw1Yubjh
LwIf7pQ4tjTTEUtNMm3wwEgYDIy5nDiw0n9zVyuME1a+sOBCUYGP5gk1RnQ/lEPRclkbMKiwtF9v
vdV8HalJrV1HVaGDysSSRoGGSea0a8NHQE6kTrCzUuAPhNO2ntS3A+wOFU1p4/i5s9k/KBzsCVyY
n9coFRIG6DDrnsWcrk6/t/onX4Fl32CvYovHcmTArHfIz/1uFEc66wfMH/1avRDojrSAsTXrTQCi
LZNBGNmcK76auOQepwS3Z3Svau4rjGFBJFu4temjtgjxMVzhtRcyYhrH3KoLKYGOhrD9XM9LM9Wt
8/aF++Rrl8MC5Rx3EFFrO45GkzCADXBhCPOe4X2fDzaxfuRy+s20nlaE7JeMFDFDQOfjcrwiHXsv
x3drRdo+1JUEDbkzJQwwgtpLz6FgfM7EIFTerYOVW6Wu+J3QDNf6N1PSYU4Xg1QnnByqGbdJvTun
3M7EeODtA01JNRLnzOI5YQttAzju+XCiExEVouSn70fcBmatiwQ5zQrg8OsLMfmmJ69TK/cRlF6R
UcJVAgVL7edsCkyC4TNB8VFP3HsHG4XoR27Bd6Ox8yEO7/ARm2ZCmf8JRG2E1GRJoBl750i+NKAX
Ryu+mZziLfFV64cTSXWuWq6eysf0zr38PLts330MRJ3EQPu3/HymiYj1qFx7OVfredRMt250Chft
HRyR40GJeIfDF6F4GMB2p2UQz3c++vASgv6tnQ7ZuFLYJtd0HUZRmGGcbwYH4CpV1sHBtZL9wR7g
A9U23BfCwr6Nayb/boz+KJRIugLazq4eR4eubSL9Nc3jiOV5Oi9wPWQ364+MYAfbFZPMN1Nyax8i
f+3d7GVSymDPdvvbC8Na2XoAJJliKDskcvAHRHj8MVrqksIiFG07kf+Uorh++V3sTv43iKN1JTBn
frYe3l42RxucGfjl6DSi/L8qomyFX9xgDFFijLvoD3ZK5MFqRU/Bu4tnGHRyD+xk3UhYxk/IU5Xz
jNaPJL5fMQJTDFHtOrqzIVSAtZnZ2RZfAgeA1I09Hn2NeYwIs1BE07C+d1slOREuG5LlVIV/rmJs
JsJkYlKmRd1+QP37JuWq1E9fEIQsOurEnPpkdSczE6vOMPSZg4JSfwGaJqfGcPM+1hqHiyA8Nea8
zQy8KE59FCAvp0DbtfbxAFSmxPYwXqiaoBLuTjOCifuAVVcUJE1Cwn3FSNq5iNGn1W+Bcl2V+9YG
uKcxUdbC+DaZKoi7yYAFnuwL9qjWQs1fuULCZt44oN47S2FY8cR7pLusx+jdYZ1STQgt4aJ/WYS3
JbBGz5I/Kg0o3Zq9Yo1uCFv7emh1ZyFxYMELZdfIrElR1ZK2pXyQmmcmPsmatR/qdgJZs85yW1PM
OqoFEsVmAxYXX6eAa80CwXP10RUTgQox/Yl3eI7EW3buVnmmhuyH8NdaOZAIhZwTvvEwyS7upupl
ZMCgjTJevwPUebj+FiYHx9BSuNwxRzedXmT/+TzR+SY2X5j1lSpdLno76IOi7qOpAaDuVMAm9kTI
mksvypquWujl0KGoE++67gkNSH5yghRIS9siBhhTBaWeF/thFBcygoI1oIWlbgxxnzYbXrrsNSw2
7/lzT+G5Z3woJaBce6HwdmHrK2Fht6irqd/a622n99NLbaTYnLLTTmK9GghvC97fg/EmJj7Y2XGx
jtl3GUect34c1UTBMYR4iaQSNquHoeIl8YFKNaQTzRo2NEvq3yex/8FDgm+8O4yjwfet45pDCuZO
p5yRCNTaZfdsId9ge5oQ7UxQiQcucUQwX8jrgf605Hnmfg+tU8xEsx/IKWdSEatvg3ASv6ligkO0
ghY2RQvfNpXi/Pvlu0U7vRQleI4wuhy3eGkdZsrehMwHszasgOB9q8UD8z2eKzgu3yKc7kaHESf8
OqHszwv0pMuRnq5IaYRJ7b7g66jgL0rGo4WMPvFjYhrJ0KaX0c975HIiV9pXHiLjgsVdTn3YzYHZ
wALSiV0+ocGsegPxxsr4zJTDxGWPYUaSG/WwITqUWtH85qUywEOSLS4pByjkghgZ6PhHlPFD2JhM
7FobphdXF1VmlGqzxR74caM9+fqliEc/z4EoiK3Qa1Dw8iEH5YyBi8wv9hHC0Tg+QxqiXvODDnHV
7BXm+NZS+mlWOgdSYv8NwrwmqV6YKY2rZm+WTMKm3/psYm2awdXCYsBbW1mXQh9y3fNBhEMbR8IZ
UBFXmZw8VPKrsIlwOqoR2rCAZtV6C8PE1ff/qQhUJD6O6Pn1iixUWPqP9xVzaPrV42mJiDhGOJs+
Z0Npetaw2oYbwKltm8/CKrlEm3vO2qu47+zIqjTtbCD3OvGpAmYHZYFqT2mNPCgmy/aUf/MMKJc8
q/m0CWpKC1b0U3mnq5q7uxvQCjtGpR6Sa5aNePAmD2aZUehr20lLzhwDOfT2sU3skgREKBH+osa0
r+hrYVPomftSr4/7bjWI+fcOErNoIdzqrLOWSxTm0nZ9e/+4ZnFHiclp7Fyqx1eFlZRwmm/Kl7ct
DoWn4ltGn1GQNPkQOMKjBT35mBJLy5WGsYINyginULLcEzbU0O9h0t6HPa5+1bvpm3ieZkoArq8p
HnuLFAV/nlvJ4ToW+aLH1yaAm3IxPKTV4apEaW/zFJlhp9cK3SnbmpQWLXbMV21xZFroFAsvv04q
WzxWfe1lCf0D6sRi70ZKEQmzseEhVfItztgyaaU/XkWDn4suPgCDdf/cESbSjI6cJt63i1sAKmoD
eRaxV+xIe9HeYCmZUpdcVUW3wdqlWu8FqF1EBwXaW+SdMUR0q+j7qDarLXFa9wjrnM10DVbNEQfM
WrQQUBpvHvguDX+lchDfKeLGKjF+GkyRweXgTc82ZJ44sBg2/0+axYmqVqygHScuwg4su9BCte5X
DI98x70Vd8UXoTOHjEUd6t1GFcmXcjn+GG+XDu954gP7MxPCWlMkDIoPQOoHj+mMT+gxJt0jEQZ4
ZslGD0Dctbw5/lnecKOI9NoaEvq6uUZ3l0ChigFJuLZB5gl4sTI6IrqtlW0lDbLFlFeVbPoaqMKQ
k0MxKcwvAhXuXPUv4hnu3wG+A+C8lPe1FiM12mptrcQAZsbobb/hADG1TKuTpk/7PGqXR1PoNmkv
j7j27UtnpE65H8Y55B11v+JI78TqNrQyGVM7+/pYWYXt+CByBON+KY0sE/ja0pH0JYha1q6f54pL
bommLx6WU2YZQE5Um3npw5ePCFKJYC99MwlXqemcQXqJ0egVthF6IdRsUcvAZZiCDL3FWpsAp7o4
2fduTctenO50TF18ScY0Qo7TVTA0wtCWp9wlpKNcBlc4AF249enSEvFiDx80DFB/nh7G2E3C8ojH
ShpZ5nkjnqwTXoCeQeHVguC2GCzMIejFFW/AeB0lN/8zVhnopT8B1wjihIKhEY/pCpYdm0GSWRtI
dQPZemwmU49UT+Us85PxYz+2Eub0MMOUpV5hHYA9X7QguT27BWqcidpKWEct5cTAzNIHzCOqqvNS
YuX/GHsE4X22c0eQ6sV7PF/WAx6+80+xRBUYU0OnsrulZnohHPwIGya+wnfcIhXPBT3+EHi59JKh
OUG1997u2GBY2cFgDu8sWTY7O0THR0Vs6WCgE04sjSyXp5denz3bzkPMnXNecoTLB6wXdhuWf8B/
7SxTzd72E42P4rPzPLfvgaLnjxlU/tJtk3HLvTkx9CmTjfku2NEoCg70qjlbbXnmeKAZjVjTnH4s
TK0N04Gck1r9T+u4cMwLyFxexQ+KG2+1JqMO19gk198NemVAzybsDemUcH997khgfGs1jhOoIVWK
aqOxHVhQuCCuUPP3tlPlbM9gLs3hm7IEbsx25ahXZkzTZcaoo2XVfTnl5Egyh4I//76VTpRryiku
oHyU4xI7SIkFgfNNuQDFam2K2gb0pD0K6OsWsox/ePswhfaUVaMt1lchX7VxUCqSLbtP++Aeskli
pRMq59Ch9Sv6Z8PbC9z0Rx/1QFzC8c0ZN5XYn8wTfx6dvvWvpDOyDT1QrDx/AbCeVluw4MPzd7BL
kPtPjDj5HP6rCAfQfYbxVPPKP1fZ0zFW3YuD9G/gRd4kvRtnyPTLZaAsbhu10yRl7wRqBLU3lAjU
FyRNApoWPfJIR6bll5fJjAWmkCgziDcb9pDhDSFLIVtBH3tVIAFVP+/p9FAfjuG2Y/z6+QE/FLn3
pRN2FtLo6EUFgc7XJtU2M+Bmi33Ag129jHy1tIuntW2Ujq1dfAE2MLO0pYuBD078eFgeb7lzEUaR
jALAS87Yzr85zSDd9RC9RWuDFxjoYtx4Uw4+gThO02MNnzUIY7qW6K+3VmG5T1tbOhcEBXok24l4
4WFXSAIE77r69BTa8kl7DfjciZkodYEs+eFURnfbYGO5q4R0hThBYMNjYPKYUuJ/S88WAWfd9fbS
Hw3TjUtZLH35wmR8nzskJ1jroayCJtoRR844MefZB5Popgo7RByatXvEhFm6suc3fKuPGDn8NXoL
u5uxXBYgv8maVOiwrSH4xqlhDNnRxoUSujK6P7DdyoCXB0xi6DVHZPZTG9/Hl/ehgfIPv9fvRCal
5yoaVJ57ATfmqEQhpF7ynpyx6Mb4J7dKj/p01jQiMiAkT12Taezw4keHvk2Fw79NDKBE30PeFdDL
xpHhqrY2TUViwDvJg5ErQEqdlR8m80ZUIzk9w211gnVFod60MLrYtauKW4fQcjaEg8YEuhuB6f8m
2X4bc6heaajdp2S9Fc6/Yk0OrjpojzykSNrW481LqHC7r5xyY+5lcMpRMWW6tjMjqLwKqGVI1Jx1
zI/DKus2UWu5MicS5baN1Q6T4c1VYaOCBqTOcndhjbVX3vpB+QIFMY4bAlgviJyr40M7iUH0nrnB
YMwmD6sgz+iVndH1ifOu8bOgNBLrgwVB1T3JapZ8D1ma9B5Fx2zyExtngV8VorLh4X07vUGlaHI5
MsKZuYOh2vO+b0oOF/iKyI0PRNuyjsSOWO0f7Xdl1i/GUWmGCaaEFvAIEVo7NuHMx3neD3eqhnzC
bVSjkU5M0+wNTHiFKFnuoFhHizMWxUGfUx7IMdfhJpcSSJbAahO0sSZ7WRrlGIKvjHKpj6/yvmY3
RIBp5wQEIqH+34tJzvwZze95+s3DZFdwXhqUaKJj2BqmPw2n21+uIGhrBjOveiT/cF3rIGs5eW1p
1okwzSHuxZDX3fC49U5u+48SDiWn9pFFcZ6bNxOlm/bZsAcUHtCykRppYhyVeMioAVPRr8nYqQ2K
/dJP+qlrZka4YFNCb/i/kIpyFiQtL3YsPDqCysHj3UKB17MLy/8Gogh0hlxfoJzVoP8kGVaZcPid
NbIxc5L4RujtqkZfo0arGWUEJZiBYusCFKeoDlsjKifIlieq61DK7ZwxpHPcf9Ziz/WzqwQuaYD5
3+fdE6LqgMuItA/bnn7TUMOIOStjVEMy4ARILU3ESVqq6+jyapdk5KxqzvksMZVew8/g+XpS7wuJ
mG3SeTwLsgrTkkVWmCxRiTfNd0kzoEUsU4g4vlTy4cw1GIuX7qwIOHz1z/Dbl1+Maqk+j89rOije
n5tuilIX51rcpKFCQcPtvLE1RQEnCaVNi0r0uoq5qlNZLoLp6VGp+6veA3OgvM3+5gsL54Jy0Y46
nUjDJqp7cM/Z6WV4DRMIevBfFnSysbo+g0E3GCliri/z9PaqghzMvs9v4zQZ5um/43YAH9h5yP5A
f01H+xqFxbrDnHBPIIFvJENg5vpRRiilguPg+JXHgu7x5DuMLqSy2AjpK1BwyDcSsRd6Zq2+udpV
Vfbnragusss8fUZA8oDQ033NByqQEDORNF7ln/7joFUkWfvrAKD0csctXwaZd20U9W3HK2vz+v8F
v2/2UlbBB+rzYzbfNAbpuYEIkP0xnEu2zbich0R/7A/X6vYEX0LsrB4vQZfolSaFgSm32fC+4ibT
iwQZWtR61tZlupvNRBiBTjT5aSttbLgx33TErPOxBPxPhqZPxES/EtmXuFRTBzy/UHGRij0DVL9r
fQrY4s9Ij4C+S+5j/WEwNZ4ym2LGIEPglij7rWdeKeNshbTRHv9oOpQRiCCxG8UW0oKiTU9AEU17
bASXU4iEHqPlTAJ40vkev5x3+TjObkbIxr3vhG6zhNy0JOg3fqS9Xuw9AwjIsB7xmKtpQxS8Qdb6
RTW9bwRRRc9qqtWkzUMbASIHQa0dL1h+EJO8qxAjb1IAmoUCVcSJQkqVOQGpS3xPJb9ZlvxWdNI8
wgEipf7rGjLrdRdB5pgJMvRPQyqgdB+i3hKBO73t+h7JXuWwbZqPteLUtmdmgROyXs/lveXCDcXL
nAF1mQnLkzLvn08vfSGRtLEHyDBjG5/6YjTazAb2PxQVmB9Faw1z+clZSPCkYZ3vW3MZFpk4Cz9J
XBBTRAOA2ZY4bM8YYKVj9jYr4HuBSV+ty/XuTOb1TdEDMj3DyB9fYeNfTCoY5A/fb9RrzCdaOfnC
p1BjxfU9P+iJ+VJ0dZ1nLceNp9yHvt+eoBlUISMZc9JPeCRYn/1s0u4Or3rMo8G4s5sezbZ7ketI
Z8pKapJbT2uyiz9sQXKf7GosMl/iV7Mf9Sivgv4iwcwc2aTJJl+SE8cpumAFYIk64tFtqZiqynVr
vd31GmNKrNoqMIf6K0FUOpozWSPW1oIlVvMxeqGIXWxlNdRUqQOc6wRcocgP55t+XZZMD+3zsjZJ
7bifqbQq8i5c4Jj8w6fv0BnXVDu3jzKmkrHaOjxKstEB+o4Io85YMuYBMsnU33i22Cs77Z3fLGXC
fGYsi6+RstlpDAGgBRlKj8mWwDjbK7H2iNpPTYoaY2x3YgM03+Mb+E2doaF2rTvr/w2ebNIEqrhJ
oNzfuCBx30w9rrGWReGlswM8EBzdq8/zoDIT3UZu+/737mC33aq81F/AWoADfq97mvn/uiT7nBsQ
6XABZzNeg3W/CymV1EP/5S9Li1F5RpHdsjIkRVm3ObtwiADy1ZTOE/u7Dj6ToTH6UgacTZAVvJ/U
l/LnUX+a66+rQ27XI5d1le4uQ9Nq/5kOEOX1IAtQu+APn9gwkEHZYicVaKhA2nxE1j5LTxEgZ74h
/yGbahkDytRwiA40AQ5IPNIHk/ptxZpakCZsHYSl4mGEMl2/zmCl2NLC5eLciq5QY903XvwI/4kd
HnagJqyo2jgNTk2+5oP+9Hvu/q9ygdJD8HElZ2zH8Ij/URDO2yq0YB2iUncfRMgEfJ9I05b3LPrS
cNR3izSH9M3ktGUV2C0HccIEIjy6drrTA168CPDOQEThEzn4uFA26cz8Df4LEjPPNLI0x+R8cTHY
EEFon7oYRrW6SiGbh1sCd9LFkMOwHaoQ0qd5oVryDNhXRA2nFGrEwe5mch/Ulf193uyrWxqMgFfx
706co50UZy9k8W6fCx1l02WF42AXM2zGcARU/eVRSNrbsRefRpSmYekjwonWtPChAAlS0c6ZLzW0
F9cKCA7Zars1BnsTql1KiWj7wK1aaTaphbWuGf3acLCAtIAS12gyf8SRTxA5deZM30hiDMpxWD/o
2V9Ca2MQnt9bGcCPwr2D1/3OXNan0aRTZm4DN1QpY97oOd2J2uvivovhIc9wKYfxm+y+vPt98g+3
6BS3LqMzIIqLDqJAaXc8NnwKZ3ObbOYdPQlEKmxe20+BVQjZQq7mgj037zuf05aWsayohNNnpXB0
GpTouRv0+g1T3sjKbhjD/Rc+xraL/jqL9SM9qBmkpVR/mi0jzd9HsMzlLGnRP8DP6uX42HC2iSZR
z+SKYan4/jN6wNvTVJaAn88bwlDHajFb7BVIcluksRzeBJYazHgDIowtIcwdV/cWpI/B2AaIaSR+
mrFIgjIFWQGrDOMe1QZHrwh9Bfs7mVm1YqYKXUP8tJ19n0l8ONGB+mdA9Yh3WNM6xB9aQ8YNSQ6r
VxF4+5RsNJka3j9kgTBvi/KTalvxfs5w6SyvhE0q0iIKQ3QryHq6GJig8iiq2q7JbSH9Xjg8h7U2
KposX1WqF0biPsFibm7HD7Uojg9q2Pu7zbZLAjgkkcjhr6kvV8T05l1rkzOCJxHT4E8cjkhDhFZf
gixIRsKARNfW+AdbFxMiQkaUn4aiZefppSIAeMT6OirZgZSnQFPrXJqGy3bX0yAdNrv1IcLul/aL
EB3wAIFErlktj6FOx2RvjVsLFvBvP87jcpUvRWIFZs3ynobqXvy9zgpTWJNjNwZr8IDa8VuX3ybq
Cx3HM36Xt9sFZHcEVeYXpNVtMBQpDRc94RhqjcONBNhyBlPbYAFCge8VEeQKTBJjBdpX2Ii5OPpv
Ois0nWlRMS7s0qiqeq9L83eSrVFSmOvNZsmg4paeVAXowjy3IgZsxUDk3eTafVjx/ZIeOAoe1XW1
Pdh0P1+fffeiu/+yykUe+4KR9VNcu/PIdd2xVOTi2WFQCdnR7N5fnkbnt6mmsUPxrAR0vjSGuVQQ
GhBe6L21WLpxIKJezD821dNF+xN3AAOVS4Mc3v3bLTBp0VrShhjH4j3orpgWa3lAygjzHt1oOveS
xH90z9p5DIjf42Q0zgKDfKIWzCBPK1/U36eAkY2QSuYU38n7/wcBj4E6N5icBYL3QB1kQlWQz70w
3zTnd3rZjGvisMor3tYU32LmD3j6S9vSp1xXa/AHafostir+OYuxT6pwDKCeentlBds6XBAo1xQm
Ifo6SOKM/7OxgpuWPy+fLH76VgKbaSzzz1gSLCnuIP7uR/UBkN1lKRkeE2xqbnUZUA4hHtWiquQ4
3A8xNtrWKurtXXW/k7g/QZ8IfaH6bnlwkA3WHwf5IGHGAETeajTefI8p6axUSOXp8Yi8HaCxTKIH
+Sr/bbPZquSXkN/gwfYHZhKrAx+kQhOx7jOEGeLbh6LDKCZaXPFigEbsRssVeC8LkMNYgrHQui9X
LeOJvGFS8WRIITxk1fkUwI9aS6mVpoyVeP930u9eN+XiMiQeqPj+kkUzw1chtWSvi4IGODF2RKvh
5vrmfuT6V/lTLUyoDu2SikLvtwJ63Z2GplOImW0gNkasdF+3lJ+YphkKIJh8IovbIot7gvPsNwnt
VRwpqx5FNwLgjQQ7IMvMkTHzy8dQ2uKfeKpVKzxPiB4jmXjAIS/MF2aK5viROouoed9PAhPIeT8f
KjBwPTwCEkJ7QSk8OOq01C9fKZgji+5TDSNebG8zyxe+m/tm3uCWDam5PJ6gh2IMaNa1R7+rbHlV
W0EpF0sk1Evz1k1Hafb7lKesSapcHgQRdRqe00XVA+aZtvzboOiQV7RC62RJu9MSuq4xlFSsAvOl
aCFeG0rR7pHHVJTYJcBBQuOkL5ShohJ1ZqhboNPL5xOn3qJjgmKuq4eUURKzFI7D5TGSAKXniv4V
fnCvKEfob7nr+7ziWZ3iirhwJ8fe0VmgCxSYcwkc/y0YG9EiBucegQGd7ll3FuMdPvswdg5Lgudh
gJGLSzVtQ7udkwwiDQvSTwS8AsWX+ejeSw6jTTFTP0fNgiRLSH4nmr8xvwyFJ/1XnVDIorr7X5TB
7cIO65gEQAzYfSKX+E65uJ44af3zdO5o/AdyIBXQzhDzlS6NMbecFdqBGXNHnQyDGJE4AOT46ETz
Ccj/y1WLXsS9enONkSvu3X7RwCwGa5KT9jbin6eg33qcwEMeb4MNFJe47itCiP+NvrQn6tgyhzQo
jvG6dELbzd0LEI5MDD8cSzMj9uniz1XQ6+bV8LbQ9r84v8pwSO4P7KmjuqGofgP33U438bG+fzBd
f9vXQtJ6i6odeQi+5SuiRl8SDqYt6PrJPZlyahqnavm2/QdbI986uKnZNo3RNVmJRFOLwVrRz7qL
6Vi3SfNcSw7griJSd2g9CBvDesuDWhAvSywEEXYJFY5twyqIdvk3T+dQ806EtHghUKz7E6ymvwy5
wMZA+34mKwXZ/fLKvXoDJqHP8WWXkWXyZqSoB9X+6m0ncgf/woSkmOKNTtI7SF+zm2JZXUkguO8Q
I5p8xGP+8MpiH1s/6b4fY/9rJxFgBai4x8vo/ERdnoXNAVTUJKsedvLc1fxteJabwuwmbLFu/OG7
/JCIYERW4kEDqjtQuQnQA5ZvBjg3Bp1zJu11rb3WljHtFMEqfPqrMCqe+xp0vhI4LrivFSGvU5Al
PS+mNomUh77pW0gAlYCvUottSXy0xA4NEy2q6ZWHRMZgMd+pHq2n6L/xmvQzOx29HEweNEE5wwMj
0saEfPWVBuFFn/HdLw3Itn5UAiS0738ff+5pfeR17W75D+bGIzA1LZvL2eXox7dPdRw1S1vCjp/z
sOs4TPUFQgRC62r495YdAoZaiFJ+R6EprR3e9KSBpsF4cVny4Vrre8GkVVryEkVP/MM5odXMtH5S
Faxe72CNb3BpZQjPpWRvtClPSFc1LAu88YL8on+bwcSqzV+LqAYz7pn6a23ElnXUL9lYdd9B/QiW
5YVhjKQ7dCc1RbYXfd2Ms2ynhVI3GUwkZ6Of31WmDlWYPS7en2wTA7sPwQWDMdSackMA6vUjQhPk
PNXWlMRodwnUjGuN7SZaLZchBcu6BDokvmSNsPGq/Hvn9KmDrnAj13OO2nAgDrtpFBHNN8cOZthW
pa5YIJfnu3FnPGiLEU54iEHTw0gd/079jAuX9r2GHd2oLk3NYhrAB5kKD/vRVh+wLEQjHRiTosy2
r3ilSJeV1JHcu+ukv8mZoofCGVrvwidDjuuQp2c7Y6/cb6oAYX2/tqBEXwLY/chA+2OWPtWkS1RB
n9I8VROerNljWT40XyT/heT7UrKQoDdS3CiLQ3poglHEaUU9EzN1bKd+Dgl/VdWABDbeaWP74EI9
iGIzMmXIGVCDd4LwLqxG+WyE/WzndL11AXPeuOt/772RUBlIslGya3sIKK1QDw05cepmdqS+nmk+
OhNqiZV74N0qVnFGqR0GctCeF78VKuWn1KrNouJYSyvXv/vRXWqIrKju7/Zbp1aMPybi72HWRJoP
nzhl2la5difjYvHeSHGIUaa8t3bQZkktLuRWnRn0A8likFLc0WCbKVlIXiPbXJcuhpbMLH2uSkFg
oxGr/CreD4LAhrQhZzYKKC0C8Jvscprr3y3xMLMChcII+yOpLDR8okAIMAFNVsEYfugrmtYcf0kk
ZtWrcEtfKDsVRR+bhCwPrTqsFiw2mjRa635cXoaTKeyIj9sNhGl4y5oxNAZ6rvIvtt3uoIhcJqIP
PY1wFUYiUjP2abXuXFIemTMx++UBT+XX0oUIyRYKL26V+SjV+eWq7jvhnDudNcHezMqCN3m42xg0
JIi1ccVN7YEJNtdzXM2/dnMdx7u9PlpYO6IGS8snqzwEFpkuq6iF3A76A0xZpedBT+zfECCH8W8N
uYUMd4ysn1VDc3832MjcH5w16Ma42pwpcNCouTH/kXpsHMFzmNdD0ieF5n+KYRE8DwZkmm4j+XrW
aLRVcQIuiUUxNeuuptspXm1kyCvzBvmLOkfoG6+KOntm7OE8mk139+NX4yboMWmwc73xRoGH2yp7
f55GV8ZLgN+xZYxxbLWgBzRXnEj+PESF3Hb+U0sEl2hNgZ1Ew9S1MN3ed/kh2/s6dGXkorQwxcJq
0nIvUYRPdO0qUXjovUYp2iylI4VO6PpV/fMVIjPLpMdjcoxnVC6mt2gmgvRvF2bNjCLr6+x8FFty
DQ+tmQZoNVT1+NSf0rkijfCl999qWnMWZfnS20qMKY1hhTTih+i5jOZBnaCOCw029HpK2sGiBNX0
qhVmQHVRCkBh57OSMv6rjN26kyvzcu1qcnXZhCJn4AwiC/18MSY2lIt6BgtmvK388nhS6yAXp6ox
iH2lhPVFBx5WydlUtkccaoGapavwJipFIPCxuDBHCH0HCkx9JfHUMKgWsQNpJeTOBDOBleY+LYBV
S46kFwaYyEV0PxSQNGNEtQiVAndXo9fXmNLVdps5ZM4PhxFAsSRmp+6ix+ohGFpUzFqsgrclB81G
p3pxupC28G6NZ45xWhJRV9ajijSW937hTcSUTrVwMB/chlv5/AgSW7yiuqiYY69vgCFXV2DSMiF0
lZlztRWRa1rg2LRP15cKqTRy7QLfnb4QLPKAn2QCae+3JK4sbP0femmBpius+V1AyqiZcZS2cc4D
amC/8kSbauF/rYB+aXIdrLYUaEyudfqQ09bIMbvir9KEDYqL1POYO8SspAJKeppfGgx9/TA9Tsb5
7q9SiKeY8CJyVeegYfQ9Y/8luVxDtqp7t23rxPS+QSg1rntfFaEsHIWBAVhfh8WE2VOd2UYGiWEd
6pPQUHK9cqD6C3DOHCtt2gUrQjklfYL9rYMSK0Agt0FMJJzsCpBHVFyv9mVg1QEp8MFgWK/5NTuT
xAXH7Sjn7JsxEtzxUeqtztW0Arf2z8UQwIJnbQE9aKgKLU8EmoAdOXqlMsv7ZdThP6kS6TamTonu
eeKgoMkjh44NgYfL2AuoYKUBwCN/ZXSpVnlUcO+Fahe5/FQQWaUlLWVZjPFvBlbSee5qa+JEyWrO
CBd3xAqUrdHRwXYMJY+GW5w+WPfcgRPVQDlakEu8jfAG+lSeXfAXlOEhi4URkDFDa2HSIcBqXPjT
aU0xaqGy+NnsVWMMQsbadiYMYwEcP1IyJQCnnqgf+EaEKPgEnlIi7cQ4it19NfShifp97nqRlrJz
qkrC8QNI4AWCSSUJP5E1ToAkd8P4dNfKQLo5c98AiHxizXXIxgA7y69S/mVITXZH6o+MElnotdhv
ZyLck61LDY6LlYUt0nzMX5yFw+qZeiZazmrHGZ9MnQmhMiepDo9VnF6Pz3h4VUjGvWaBOXM0TYcq
/BsmDrZPkBatDoedmCXtkQ61ZLNnQSJ9yZ3A10qbSnbUSoDlhcu9O4nBbznRcQaQ2JQPRrY/tYyY
QutzOjk4VjLs4EErP5kyFLU8orefjhiHjapD8N+qAtRdfCw1Ukazy/VxyOVE4pQVHniioFeJpjoT
5Jl2kIngXtpAMyDQcZSQf71eJ22iXFsrZLO3fc9RfnQn8e+6Ol4t0K2bY7ro/sc39YUPsiDC68H0
APB8+3HCXb+KI0/wzxLQ44HDVqchnQH7KslvF05fPIue2iFsQaRwVUF37ILBtw+Y2hOVkbBPAW/3
G+rPB2F165BCKZGM1QKitIEpr+kOJXCDRisTb08HVtGEUm9+7Cd/99zuk8WoheINFh7mF1XvfL9t
v8PmnvVuO9dt7Qw5JEE/xC0+AZarrBraeIQeGB2PZlgI/X+5fuPPeWaGzyKBJcNiRoMnLNhv+vxZ
0ha50YzJV+Figs497XyyPta/LozAk5a8tL2M++tZQhJ6xfrx/ZFE+diwR38gm+BqHGl3tfnCXrEZ
c6QVE3Fw1/AsNPq+Qw7kGsUK2axluALEW99FNze41sSDPEGe2ebGSVIAWeBJSp55x57Ffun9f/xW
5zwnct9uERQnbVbpmsXKvJ+adIhtrbrahCZSGBUNWH2aFJNyi1g5YNvQjYb1grLgIq9YqvU7zyyF
2CJiebsNiAOlWa5n4byTzIkgYRgm0NdbRGXf77vGiqRqGqID0rntgJcPOxbjFCjtMi7EIR331g2W
XnQ2Sj4Gi1agw6yMeR1CWukOjwHt1Zs6owhh5wnyHabnonB2Pdbj2O3NYt3XwGS65dBRCUpQimrj
1O7t2kQ0/bCUEmkUcdpGp6hHmmGWPbI0MdKAsDryE2gHfwCsTHfB5fTisdcE5dWVUg2QCoVRnMwb
WiDBl49KSnCVkP8Du3g92QF+ynhIg1zE1ku+9cEaakmw6DQgFPbQKvFZisPv2mky3FoNcWmop0kY
leb2uo+cS6ezLsFyaqFMH6nBcehm9/VUFuFsjmAggAf7vIUM/jQYcvqIvcGO5OFkke+/3KMpW23p
6QvuEYvd04grEIwMXQSTNmWNHvZ15+99dgvRG5sPY0NKS+y7MzZW3JzVaitgESkR5BB3pPiAjAc0
lwbRIPXv10+ikKVpA3S6eoAsGh5oPce5Y8BzHlXiCtf0Avag29rhvxEuyhsldslKQwgwfB/LuCpM
TXLpKcbfwSQ2WhO75kkZa727VlCmK8oWvVMuKGHdr/yda1/IHcGc7UAq6VJGhN0r3vT6MjcSzJ6V
ZC4Hn95Ack+KDK6sP0+wPjb1bvRmu4+WiUdD/997aOXXQ8pTiOSybaUeeeFz2Bj+OwM8B7yatSTp
yzSfjA7MDatepaAUXS4p/7X3sdgIWS4x58UNeQtDtKDIAlRmaeA56QQGMs933tC2NXY0W1tgN811
V+Pby3q9oBhDUqMfHbImPT14JAwZ7vCImjqN3kNp/ZR/+nDjQCJ9ev/4p6MSKZ9GsLhEAwhVinc9
DpfnG6A75BkccXrGqVafw8dlq4W3qtQaW9LP3kui39Wp/S31kiuBsJACLI4soumU2Yv73szuY4ZA
dq8gpVj0Lb+/KULYqbV2tF/EIg51FAMmhckyOLfspK8qBe97VvDKVloXY0Wja/F+ex5jXA3+V0Pa
W8GImDGnGE9dZtCypcFWjD2mfy9aO4JfYvHsMkiYiUT5LpcPJ6UdH75QUCGOC0bXnq4BBaftpVTt
bS2LRfYJmOIVUaEQHrw+2T12gu8OqtkCn50OvV8WgEBrsE0eZZPdt5KP3ZQaBPgoWC+PPs8iUZzI
Mcuxq36VO6xmf3qIZCdRfWzduLCXIepGtiE6Vr4ml6JR8e10ZfgtujvQHAIVZZ139r7wizComoaD
niMo/vxAFsjRzadmbKPUlaTj7h1pb68Xy8edLL90cmYv4G0yl7+Yn5jWLtSmCxUHDmwyqJCSigUO
ji+g+Au9MZF96jC+lHH6q6KrGnr1juVPpCIbqxvpRHoU9fU3fC8sXzAvX8vXOt5B29+h1bxqIWOs
gJNQ4iiMvp5fXyYLv4DF7dKPy1aoCxsSn/ToLy8atmnObJLfA/WYf0oGAvk8YADHiKUQs/E4V8pL
zY82t0qaEoqYPT1GUjRNGvNFJc4eId/pPmDoCdFX1PV7wBp/H4gfCD/GXv5WjMeSwm+e3FgN0vCH
8FTEL3d+r7D/C8ehWjmUEkDLqd/pLzMOcscPbsJZoLCQ4mpG1XkE2cbN2AOGZ3MmEcFCVvBxAibJ
TsXDUUzHFpP87EdQrK9OWWHVHqo1hDJpuYh6x2H4FvXWxhsaUS+rc+plyMtQCq9gJCcMaHlaiUpa
1Mz0hOgjPN+YBsqfWZxyl99rp6lbtT48ZqRvNGah5G9IJ+i9VB53O09Yd4b/YezKLm8cfrFXRDCq
5DXcCp0yvYeG+KZdVB2o+Om5gOSiQqX2mee70HaWsgenDF234sGoKP9M4/53a7b+LgAiC0BONxU3
3F51fS3SzN4fL7/bmlTimaIaZKDQiYm6U89yjGIOpDublabpifbqecfxNJ6m36/pk0Ap10tHYi3H
4p1D/0qVgYD3EwArIxwzgzbGdGXvbxLpRacZ30BLDb+uzTRlx07vyGnQHPZ9RMbVN59FuHbuGyo3
P2J7OMIkRry9+yzN/y/WUOtYdnlq8axoY3NZ2heK4JfI3NV7fz8KdejylsBiV46bE/KazICjN7pL
09Z8mUYojP+76HXCFu/DBNZelnqLfuFuGPqcHRdVCx0stHOfODth2ttNRAcc6kx3gogJRgpcZW8s
xAhXqcPwA+z96MdaRq2oSUd45Gv0sEGaW+Aadh+W4Z0YdQp2Ihb18XeO6MrOdN8lq9TXfoZQwwrT
SexT1S/Pdz+6goGM6flOW5wk3PO/7xTPHVw6IG2ozcWshnyDIZjEytqur1igZ68Hj8gvZksXjTvS
+zrLxJuA7LlKwI45d5KnOD20wIAiMadYUb8Ss7rct8Mee1Bza6GhWzAL5bliOo4uH0ig8GKvbaY0
3gxMvjLWs+LWPMeD01gcSeMMDgFDJphNqMHv8NlFVmbCabilXHS1+k31O/etd8qGN5seWap4od56
V72sYmk0a0KKis6EDpx27XadFRXCHLcCXhj5p5cgdS9eitH/fhe955z9q8n2WRlvP3/tNvhlAXVX
nCVaHEKOaDPIGz0aCkZZ1MCD1VA3QmJY/CPaUE+A9GYs3Tm5JYxW3hHE45tJnFrIYLFnnf9vjLP3
+Uzn+00Jy7JyXL4RbIWyw0Yn4WudXqTGTqSPiFyzbeV80jgqj0pfpWm87CQk61JtdaEtISnB5YdN
ryUcduBIr/qZ7R2w31UCUmOwXMAbq8KvJdVTV3XuMOl5bAtYlZqHVbPWqfJPg7MFL/8XcJBABLV5
QXf/g9CTDodx79y9Wc5OhvvylOnRdO0wLOrzem+WTkjXKfUynloMFfb09GeG3zCo4ZoC6pefShYx
PQZRacI0zLp6OBdywPacrFQlPa7crvU300n0bfcrjy1ZrbH9EwF2SKars6QXYrARUJWRKFI6aAUH
1TWU0BTs8oMZVeZl7jhPZBIgNxdMgznsTvzkMDZv4OjmRO0LiP9Jbv7MGBeo4bjW2JhACeSTjgl3
0oJauaw2tMrj8tUNiQPyifKW7WgpJfKw4A9HVpS/6vo07R5vVAU2fA4CXc+jBJ/hTntpKi9ZrjLe
9ahQ/gQ4whlf6o2pBmdDdCCvPm5EhVaOaluRtMc5QkwkosqXqffkpHvJMg4R43RgZgxAXoZdUnqb
WsS1ERwrrsxzA31BOWTjqtVJb82Iez5GK+3WwWsDyB4vlpvPwtgcANhzcA3Cp86y4Byrpu+Rbr2L
CaZR3tyC9uyVHIxLjzYphQQ+RttAiVDzPjbLiWrA45K6+tHh291TvfL3rVd5UBZttBt+UoFe6hnp
/mzAsPMoEEmA4+EVDrqE0TLx4r5WKRRCxyqmYW8+s6Tb7sNnGlEXE6l2r9TWXlbu5PN6OAJJU1WD
Wq9n4utZXo0YjY9udEGeBZBtFTLpH9jJ7cLoFALRKO6yuCFWZnJmVn/BroLmAIKqzCz3JHM2PGIT
GoXrfCHoUZXrkGgEALb7ZXvXM+BuVrh+VTLUESZc2mVmZcr4pwV+9VjE7mdNgRB517v2nyeSUBqV
QbLywjf1MzuqX8l/kvUmvbV8swTNfdpYnkrVMYxVxppUYsvDk/3UYTWt+bPW0ZDhdsO5eQBj1eq8
3qBialA+h6uDy0pWRWfi7kp0EwUXG4DwdrB7Py2GfuAVBieoGk+vIiFz8nk/Qu4rbt7mcBPPnXz8
ZOg9o6rG1JZkQJ33tJfabIeyWmtWuWtfjYDeC1lN7q5xTWYFPbz0qKbL8IQYtxQwOIXW4o2FPQ22
gRFOEu60pqn4fUnnx9oZR7VtbmqKEUKmc4DyqgeKTTSxu1QMDOP3WSUjMQdQa7/ldIEGd+XrTYPG
VeOyQYzxoBS8WofRxNJTrzHL4U0c8gBldG4qJTuaMu07ocg2bh5TUUgGviX+a/iLaOUqXCsC0REF
8cXoyQViqoTQx0l5nuwVpp2DFNn5JtwbgX4rTP5j7LlYcyAs1oN0lFalPNWgwC58fT2l8Wnj5BrJ
orE3HT/st4bURQtv/NuMuLO3qwYOAnbQGzS4olZ3UUo9ouI10jv5LiqaGrARczmU1a1aPSrmY925
X/Cpwn4qACYsOrR9zla2SYztnI3EhlPNOF+jyrilDwqR/jhrUXm5MMvyAA2X7y0tMPM1c0BS9trV
FFIbQjst+yox60C7fJTB+7aX/17B7Z+4/x/S24j5V7Yf6GuAVCZRP/MQNDDwdzWzzxXrWYjnSBNK
ZUjInAP4oPMlJyWSpns16yPXFgyLV/zEFAKv4P5ILmlgMAB/98/XzFxFQEIy8y27Eu/ckdbJtuIs
nb6AExCzRv1i/x89bo/novL2q8lG9ihjjTgncv3K0lPMTT2XQ9GLpgKCFzlLPAfg8TFheeGYHBpv
ur7oyCDY9EivXZoWRZJZ4rS2T649+MI4qLp8fvF/W3X6AaeoA4/aD7Mpk144zfkI/lKYdm8iPiPA
g52Dd04Nxme4SfpGGPNi773elgE1uh9AglxaPe2fVDFf7tVckIfv1/iMSPlsaXKnR32VrncvW/d3
eNP0pkb0aNqMLrLwWFc6Wc1txP4zoFDRkn79FSganyfBgr7T9iKjHj8ZKHD/KUStoccE9YqR+v9Y
HLBGweRCgRQxChz8bcnMu4/uszNP1BpB/ivua5DgkAo4zP6MT1MmweSU+z6EJ0x4aNjn5L4/qiia
akC/1wqiEbBU+a2x3F/Ld7XxwQgiRr1edF9Zbq2bqL2oroPshBWPNwdqyuv4/yYJZG9j6zJlAIor
7PEDQXYDORqtJ3ZFYPfO0svUhP5jWNRDsZjcC6aZF6ZI1MCRm5jARz8rRs0NHaaAymq13rzU5IIb
D8g1ZLCQJkCfGdlK39RMy1gvP2JhAyo8LJJEB5mpmSdJ1E1ym1pPU/oUKJkNA44PXABnn2v6Ban1
Rlnf94rBubTBfvfwV9gz38ThxY1iMrE00jnMWmqbNZDwS+1+fjCHsxyCk8JU3Ruj6ETuVKynlwGL
lSGMm3bW4uTgpjEcaRush5zXzFZ6kigutW701T3L+Udq203QUTvtLkPYWetdvKtGig8uoFYEFrWz
lj1FRCLOevDS/dBltMW0gauLNyGJ+6M0hzNNYfqtyrXemSHCniULjj/Z7GHmNyVJt3gkuUWGGYM9
JeDt9/8BiCrjba306YfyyN9Ehwn1ktSLAqbMRXjLckzNyzLvHbH4jN7m5fOgyRtAi5AdozWHuip9
CV5pVDEEMYBKXukhKVmCUBxWd6/xoQ+votYlJyuCzTbwj707EegjkxVQLli0FtyQqnRtSk6HWd8j
mXmZsMDLr/OPuRovaAWj1kxutcUA6AS1lieutOkQt26ClPN/Y5+yrveqFQEPIS/7aYAfHk+zHi/W
/xmTssWy1lpmc2Ou5OgPsLO361ZQkS07RgpbKXHOIMzN4hJGmTPFYgx/h+aARvY1dfuUao05Ze9B
3r5lfh6GeQCWFqtc0aro1qveLaLeU83nqywk9n2JaizyPNPjEyj2z/McxIh/EH51Uv3vbzoZeBye
ZXp7/CmcV1610yhyBRLJcpkrvMZ9QqVBQ73hLltc9J1ndQZ/xPopZn3V/2NK8wBo4NT81TQcl7qT
O2Amo5Ohp838kttdFns3MKgXk+DYQgZMaLAPhU0Uru2e5t9yM5D6JEslYsbm5qXsxRg//gZN1MeR
1VZFXJMn9w4wqgNpU7bblDJ3OKhMBLnsGSqt3XDXK6Ci2aeMGPQ+8h0Jo3f5VolDoqiGUesxnXtd
TOjOFCGUjMVHCtSs7atASeiP63HQ1iYqonUNyEPzhgJvia1O05kLGui5kQxoY5zEdVksvZPEP+DQ
SGEShEUf7lGsEdbPxEbh7jQPkz+L+gPhg0rWUWxpac/gwIT34OfuSBlBm+P4OtnYUYKFwb1yN7qb
3YgOX3IbNbuiobA1mw3fPUWBK7yl6w6O7AGaHmEITT54+un9rI38AbLIUFceomfFbRtjSZbYfOeN
1rpon9xl5JfSzica1WpTtUvKsBfqX3bdOvMU0Ygos2gYlq6lW0yxJTwTby8SCqCGUoZARBUyYiya
VWu60I0mKrvRE52W32osFX6fIDzjTWAQWjowUs4GLzgA+m1xgHZoc9h/+WYfFm8ZWwtVepW0y7Ef
NMQ1dIdF0T3ZOaADwnXmesuQOdeYMtj89D8CfSkeWaQDJGuAgzUb61q4qGQcrUtnvyYZfnqJ/ZfL
+X4NmIjtI8cemc12lWiUVr+yrz0zR+/Dn3+Q/bMdYI3OLFfV8+CueW2ANgfPdLgcdFb++n2/htpu
/qGx5EKkJoZo/T3Mdpjy4XPaUc28R9D/S1pkPFzS9g2QEEO4kpLsGLynQJcpILLlqMFEf+CILwRb
guzjxAnDrbLks+tvgWnp4eHmOueclFGYPmPGPgIVxlFpSZgvuqkRh8++wP8PclHUdNLlCwxD2D5v
vuVwaFJLybdfOMapmc0Sp8DsdwVDnFx8xbBlcjkVo689TlqES5z01pcKutVUYdCWurDFwsWNKbDR
gBOWS7++PRtpw2KcHe9JVcU3FQMyppneAFgQqPQ7xRern44aK+kkThx5SPqvNsq1Xwxv31iB7c/+
7reNM036x7dISvD8jv+hFxajEiPHZSQS2HeecD1gRrAm3628Fd9AOXKWuouEumVA/+MasjIBBJ3c
sIJHOFgzkMQCdeXXRgtt6afRFRwzZj1ehdar7f87YFpvImX57hsVfXCBRW9bS9R0jz0NnNR+8B9H
i9rQD3J/itz6mOQRP3KxAT/s96xYBnQ2UXFdz2q2gSDxgCoGeMQUnrODlKIOUyjphTPXcViY0CVT
Uspguf9UkJWUCDEEjwAraxvbywL0CELY5yhzdTL8+NFV5/6WQQKUBNfhOoetZC6NDUL1AbRDl3ys
kc6iqfET8g8rmt8AgvcWOnppLe31ITCzc6SjQrnVJMHuZ63C/MV5myvn2WuA9u8GAomhkpl0BvDk
NG7OBpQtu15ld6dZAnyAcTQNXehs7c2J4wx4yO+gxeUH+hLm8XXfSNJo9jRk12SHO0hmxesrbrsm
4R6/qYViYn2sLOgifX6ubNKQXXSw6p3x0k8+bpXV68vtXStyy5mVAirVNOAVEQkjBUpzPKY57vC2
jKSedqzGfO3zxIO9NfawyPx9/NGmSKcDnt/WZKqRjZx468CYHAjINGpvNZX4dL9Sxc/HpF/7URq5
T48Rk33qwGadQ5AP6TxBf63zkR/4cqodUlo8yqVRfyzSZTSjfH5IaY9Tw0BQhwP9KFnTP153U5jn
5vVYa5T55/i4kDzD7+8jPVtP2JCMC/CWy15mOAlRPMBvizcRYngaKR5ddj7owAwjJSCnZgMnc2nl
mgLZkWLPMbnmXHAXnd9kXNNJDs+N7+/5laI+1D/+oksDvJYt6IkPhq5RPDfSQxwGR2KBlpX/xQ0r
K4wbZGD98wT5xxMWNjRi/fNbAHNaZFRFi3CMrA3JhbGEHOOpCoeCiy7qWWKQp1OaqabrM3jNE/GS
IHdficOoE9VWt8givxTGawv/MjbVA4me3jP1mQHos2XYLt7R6jhqpXU7sLf1bX3a3dI0dkXf7mX+
xodLQLTTgyscGLmtY7XOc9ttoovbAp4e//XSFggNrMQQBzE6+owXfjz9otV1MxVDwyir3NYoCiXf
8arm2OpAQcOYadEFhXNUruG7sf2y5j91PqfVP2VDiMYeRmng6+Y8MPqd4Kvp3jgAZ2VTVeZ/QIRC
EVKui0DMOTOSkYLLx1v3SSfIULBO6B9s8KHT724Urvv9opA9IdOkO7hZSesSiL8FvIvQcw96MSeW
9vMNkOPpz0DQIwcb2i6CMIH5JSBuvsORNgXHzJQKxKxLVLQvZSWQTa8xqUoCMogwt6XlTL3nrKYX
hEN06wZuAw1UqOa99Gp0OryprsNjYhpRh4e/u0sIW5s8oXCGRh6FPp2rPzk0LK9IrZR4gWgoVhhC
O2p4LOYreuARAKSzwR0jIFyLW/WPBG5l7HHH3s4twalBRGGllhROQyAO13a9EOUK4v/l9o+G03Vf
SjHHsSJeK2N+p3Y2b+IlXc9hJnamVmcwnLiJHNTH46f2eAwPaMk+oez2LJPBuXu2GpEJ+ixK7o6G
u66/kYC3yguV/C0PMCKMccVPIC12b+kZ1wNjWHPzzHQdsud4AfMKVGj0faLyY7hYRkIc7JdsNvna
XEv8X6DX4Jdkz/AwAvVGTgpvSBQsdAi6hA+0oQNTZ2lNlOYl+f2Zz8pEOcWAyYzpea6OG4zbGnhb
dAohFl1oUho791srVqXmt1Cx3vP3izoQEyeGufi7zal7mn1VDR8wRvKj8+FWPUO3L3tsNdGsy2F/
+qK8PJGn24wCSjzQvUD8eCI4C721iz0rnuqwX2m7uNRfgRYV8X0V9IvEMhwa6oXA1jaSlwk5lUz2
XnRl8itVplmr22f/bE2UZtGupj/ee5vzddDZPxqT6WcvFIylPJPHbyDeBePklebZ9r57wbIDhb9u
fE+q13gXjM7lQt08Vu4Q6B5SM/M3KHPXN8veDln3erIddJseB2aHeuN19Ibmz+smv8bGLP8dWtj+
/blzrmuBb/bXy8NrurkI2jy30gDqPFq+a5J4/xAAXlcCeNh70IbN9x///AdoN+ZC4d55+bQlHIFS
hMGydBMUhvYsyPq92sxIga6cKy1R0EuBV0mLOxWqeCjA8ZI5YSVlvr68OsJahgOpRSy7SdWktK5W
ZXIGzEreWc4YhRB5l7eKhrxH0uOWIN4V1FAQJkE0us0GLhKbel4Rq/mbO8OGY8UFWHzvOGO9SicL
laOfRJoqx5fu502vNchFXWKKZoZSgTOWW83DegN4bJdzvjGjfXiXiKXTv/ZtAAPq+yk+NcEEfso0
8ghDRarxM6D0ih85WqQQIvD3f5QTfmQZZ2Tl0GErryVrJAkplcN1Ode+wXmbWr6YFocF7JKMthtY
ebn1cVJvz6px3VYUQ8O+ZenaYSxJj8vNzgppLZuFrkLFz4eTL78cmGpp1MyyMp0aA1K/tMBjAV/x
Gn5SpCvr6VM1i54T2w7SkCN59IY76e27uWNTld7kJJF6WZ8jlSL7AO+nfRw8x1csbkFogA2tF0EZ
U+3tWFGnJ1zYguAF0vZhdklT0aFoKSj6OMUr/QfJ3b5qRmK8RNVWL557YaEtRsZdzd7sdC11Fmu/
7GUJkL+rx5LmuXGRhCAYboXNtcgEsdyNUnfNJ6efW1ZVkqt0kOnwJn3CWszifyac9FBco6njDfHz
NSMCRZbsfhen2y2wvZukWW0l0jYlTNUtLwckF0yl7vbSwxC2ELjBGhKyP71HF8bm54LeHEiH+UzQ
EEd1aXCmEtud1MqcG7TC1cJTu75nEtKZcledqNLKppatSIpl4bnqVBO/4NARZkRVwPfXTMARNZ+k
FyUdVHyW/nVsVie5IY/IXZiY+CwwsxFne8l1F8zMZK9xWV/Rrdr+YAogNCzc8v98FrmxAzgWs4Ce
fsf0ZD6NBAxLoaolN3D7t1IsxumM3HyUtXA/CTCYggjfZ+NRWRvRzkDagVowVA4fj22rNhPNEHMy
tKrXZdNIuOQdcJwvrY31IhQQGlL37aMiFAc4Oz48POMgr796ltfevduvsFrOSCvJQeeMqw+lOR/l
w7f9LsLBXJpvqEskP290ZUK3RxWCodmcjhG68BwC5b274nHHrjXz9JtmED2HDKnsBh9s6MUdiJhN
LIxaiyPcWgACTt8XQBKPN26pbNSgRoVSh60evM5D4BCMeRTs9X/6fAPaXmhQQaiQCoIXAM4VEOXm
BlC07E6UXQBKui6+mS+P8AGmwz55S+hwSxtByxrQR1nNMLM5TGMPu+BP+g1uEMcCyrAIfCc6iP4N
5q2UVEA95x9Tyq5+XPMX9vXNKt1FjG0KwPpkJOhSMUwDfgAF2KvMFU8RYS2Zelw/Rwbh4Z/4jz1h
A/WZ7GtJh48HBn/JTwriQir4GdG66uI534PwNLqw+GU0pf2H4lk9A7mtXAIZqrpojq1LJc1fj2kR
pWuMdnLR8flb+BesDDLEov1W/eBIfPDfAH5Fx8wXMOX5Z8wBwde7rHN15x7DcFKzh9T87dgvvkjG
hXsCYN/PT/Tc6cRbmuGdTPThyDAUi2hvZrBhYNX7rFVdtRqy+0/Poi6K+jEd3iuIrqyD7ZiikO28
9htAS3nAElUj57bk/I9Q5+aJwlEjEf5BDUU+aUJzHTw20CRhebLrxl+ag2YG4FAsdGjgxfcD1VLb
jerLs0e0kWaGr1Q3253+IQQkvdTU+3IrxYLEot7BzohVY5ZT3WWNsBDRL3VITyx64sJtioYpyqp/
1mt4m5que4Mut0cVKeCVqq/lcRfrw8z36/EeSLem4BNiB1NuWKFQ3fCKD7x5jCaPMQJiHaJ1pwUg
DSyh22gzYKwgpjOeTbk0aOkFqQGd2qVPeJTHQKKOz87dFGo89oebroDphvQTqlJJAz40FIlNIPiO
iQ+umFX8iOsleFEM9NKlK+5zoi3RoSqdjTu8aUMUvgKZ+fLfo2CRRFHXLR8BHhZmqJPPjhRdtGrz
CKwQxPazAunFsEmLWqki1nLKluXN43iXiddufKl/v0XNPNgI7JX6tLYCJtwPI4WpcMujnCdsgDjE
6VxMI7ffXIbWnJO56DlN1Kfp8hUtY+edKpQOES8VVzJny0Bj7WULTqWxjTp7hfl148fzcdK45OYj
0rD047AKxGH5xMO3OD9Ge31jMbSpIkcdL83beW8vr+QgUgQG/2CWbVVaySLJr0vbDbJQhILxDxZN
Aassh+5bamxKJwdnh/rdXjA+acwykhmytyEeETaYgHiUDK+oVP9na8rxE3UOP2Y86sm5t+BQX5e4
LpYJ1e4IVUEIT7fFC2YrTV4Rjw5ZYpAzFev2YX3VZ4AxhwOkxp6XnYA8gqNNehtaqfKpzbHaqvAc
xWuRXX21jk+Yq/bADgE2z2PGjpDDnJrEZOC06GT35QBQXCUk/UMJgZZrQzggvb4VjRxqlAf2HyuZ
hJYt5sx20c0Zg8ES5eisA9/lzC+N3bwVtniNSnlb6rBfGihAELsbq6KGalY2u4Y6gK+e8/9pfiRn
XvgtMJ21NrUeKNQcM6G447zWXoPq2WifmCNetPHZTxAJ8Kg5+HDfn2jy8AF5t+hEtga/veIC8vga
nPFpAf9QBPXS/mOPAa5mjaPDQO3E2oNXXlFGiLMEVm9Mm7JT9t4ffrjogO8vNcexRSLq395+uWzv
Wg2yfG3Ov5Qz1UPCkKkyzwsgESgfqoJuj5lypcuMXU2AiBhIpdftc30LbDZmN2yRu9eWNRxA961V
8QtGKlu5nEm36tOzIVsJRbNHBZwZhB/EYOnyPk2b6VcGRrhMpaIkxscqgzlVH5a+qIPEq8lAzVNM
1STNABA9zutyWaeNf/WinvOFhwV0eW+GWzWW9LMkCgFexSwm7jlCY6yFoly+Jd0UIAB03iUgTYmf
frm0B17ElsXL1zB4ON+mgGT9/l7ttKbXwsoDfVw6c9hR3FEBIgoNaslAEXYnhcEzwbnw5axIlBui
CHNbZrsHYSK2sFGOOgpQhU2s6AsabADyF1b8UoVniecVYeiI0g8cAJXIhcdVcnb8vo82s5aAp6Ux
tGOVTJhGjhDxlsN+y7yF9JaO0hJRcMox86pUBW6UmJMlNSx4xdVLbsds4IfZITbSrV5DN+CmVRXg
vEFefYgauvSDkmAaEMR0/mZpDTSRiHvPuEbo0rojMgjxK05KaUyPCCYONOjkPlPUW0N5uRVudnmI
6yLhx87Rn6KeW5CsCY8tXKCIS6yT26v5ZVm73tXE3f0fog1Of63WJidV+wz3pm3xNXDyrcge3xXZ
8pBU91rbZ5yez9H/AtYcQxFWBkAcq2KQkRhexQUp81VItboUVU+Pzvu7BxUIPPd/ZIWao2O3jWit
WjdZnYBsCwutVbml36hJfWd+1N8LkdB9QdTLfqGhjKKRH+c4r8aOncavAi6HvY4hfBIfOcx3bI6b
7U7PW+TmsCQv8pZfR9g2hvy3o9gJLcf9KkDsKn/N5aLnXUB/mb0HI5j7CQs2eaOBAlxpJtu4NSN3
Ut8ExLzIwJl0i5aEFsfx8sWR/l+UbH4jLLojjfcvejLIaKqFXXeDPlZ5Q4wgJghiyrCTIcmvuwAr
YUUCWchgbTCHPf4YnXwzRZeDHB1rUAfPs3g6AaFT1es3Y7v7HDAgZdWD6I1mAUH2YBWPxwS7hsin
FaTuJNZhFsSbGArsOtYrrKLOZ2537atdXIgLLMTArKTF27o8/Xq+CvJ3svcwBfRBfYS6TFyajzLo
UtByGObsqazaKxwM9LwqKOhALLbAHNMTlgicM1bcAI+EUJgU46xttEVpwHroVMV6S+VVxeg+hk88
2gwadMAyMfeMAULtegh8CfKKOoVwCBxQwgImhIY6MW+9rQSMgG0mz/QSfBMZLYSnRpWSeG+lr6UJ
MXW70fDZuA2aMypZNIYkcIn8LLFA/cd/kVc+huViPC/vYepW/q7P0OjmYbR+wTiTS+9NMkitISuF
WKbiwHNdbJ4Czi1vgcNxqJ9X7yMvqY7H0pR/4Rf9ZjLy2zzVu1uueWRdQ8SLafdKsU9+eNsY7xWj
wDzX3PfCeZVhTrbbl68Jk1SejGk61XrtVQFlEsrA7gp+l6PB9Bv119TWQOLS395o/qF8OUAdEZL0
+h26eCPLynCPFWqHLBc9GYonw4PJ5FfCO3mMeGfD7KUcmvNzpwIUvPYS1LtjJAo4IIahNGfGx3rk
VphXwxffkdIfkw61YtSrKps1KoaTQZfoVrpt1KpS1TRP4gsD+kusCgPvbe4GSsl0SXqbNgmFFzBH
AddKqwyoq2S83QydT7WGho2f1ct7RcjjCGQrOHPJxGQEbJ+6AXB4kMbmct9X+3puH2wrT7KKDabW
5WTXtVBNjtsA0gnW84jEIkov1o5VpEHp/hANHAIdZSP1QpFG1bJ5chMl7M8EPRMGp2Hh1kM32oOD
7okonoxbCSn6UQfObexF5KIq0xsJm3D6r+nBaZZKnvbqTbjgD6NBSpBRlnZH6bwd7ka2qDh2NNT1
3V5ak6Uvx1CuFJlx+9CJuz6Xb2ypdY8TymnkrGvto8Jk6Z3/6tEAxwHrWJgEIa1Ap/eTJBIndDIq
oWDUaZ9YRqVjnorBLKrp4o7PRsJASbKiZzccFADtVaKitjTwv5Cr/r8268ipQQKRciMTWNiBXHtl
oEYjzDHl0F+E4u8xPFiDtv6EyqCbXKvQoCWBub8o97dnv++7nl945AdNjnDAp8wMEEZjrKU6JuiM
FyNEZVexxRDAhmzvZgwOxM+LWB/lNe52JwfYeslBHuPvFumI4w7gceKvY9B1y+RpHorhJj1LRmrV
u1Wl+MUE8EC1MAnOOC4FIQlhgksLrXSiJxeyAF0FJSYgIUUS/LZW+EfudDTLbqlyuWoYYDjwOhMn
jctCTrfnI7LXpcTCBZplu4OwA7Vo//V68i2us5sDFUsv0fC41UVgPKitDS6m3aZ7Rn3EHMwkvbfu
rbDFYHHl8oIKbLyN0L6/l4dGmqIvEicGnLm7fnMZyplzFgZAfErBDnObtac+XPWba0vBJ9Bh3b7/
wSegfCEaM08y6B9iGVLSBSzYD18211KFRpp8KQ/QF3MtoRloDPeXLNB+UaWo0R4O+1CtEflk2VQq
kwdLcIGd3vGBaMSp6uxYT6orUMp9now0U5eqqs15/e4mkFnt8xWsTq/xuKIbTVzKw/l8XjOqroeI
HWrtiWNH0m9eW9WOdo7ZmGt39MhXjRu7tc/oP0wBWdbrvhV+/IPLS8otxL3W+4dYdCOiGlySGUlp
rf6O3oiQFwgcalAE5BosvbTOO0el04cWOkmq0FvLxPEqC1Jz+kh51h6g6kGQSPupZ9pTY7EP0QIv
r3h565hLCcemR8KQTDrVs8mj6lAy5OXx/4umjmw9WlAVoNKZ+Mo6FaEtIisZ0gFwsaAOF+lb1X6S
2wTpUBwmzxcHRcqTYXZu+pj7HT5jBbFwme2FvJhqe15wbY0Nh4sVbglh+Q0kqhEpOLxi6NgwuGxa
oGjdWoGCSknbhW3lkkrsY8QrRAG46ZxSloAg84XQCqcVfHnuDU7LNk57XT3buJjeBje3pROeZA/R
OBaOMtpDd5TlTzog/Mbkqjepm/wSM3poZVuVK9xmmT0YQ1bpip7u8b1HWVxKnn3yQkjbDwUCuTja
7i+oqBMoihWvxZ2XJHkQd5i1rJR6SPkYDC0yl8iyUSolmJpRxRZC1Jwfqp1/xcGPsLSC8GPzNmO5
HVgu7xb6SbR0kx9vpX2paor9DoXHJH0gxzJbtsgYSLJrUyyWYHd1raNT+zHXtXjCMZxFkv7MWdTJ
96vUVaNEVT3XpxlAAGpUhYVhdyeXqnrYyEXbGPEfXZ9trVVnoP3H6IX0qrN/octFpQZscH2/GDnX
4OrUH4rJg/SE1ViPUoKiM30ty4pPZ8Y5zTnb8hNxFo22mfxoFpBWjrj+hXJog6Zwo6kT1KyGiNpG
rtLSKt4E9g5JROSgitk8CfFDDfh66yEyISG+EJzAwG9Y1TgvMGGsPHhC/Kt0S2QuoL8Xdbt0pMb8
0jgWIRO/NUYWwfqNj70m5FOpAAF/WJRJbD7qqnz5de70ZHz4JjcsF724pJHweAVR1np7DC/wTfcI
jqPTYoIyfjgSzwTyAqDrM5KYcEw2n3jpO2b6pC76qS42AW8Hf+roj59oIkV792j6zaVejQe8I/xD
NJiZ7K5un88GOxUbtVI6aOiZILBkD4vGdAPssUO7vKJ2nNZsDBB2M5HnAOfz2VqRdVE4sN1LcctU
iyQ9xQVxTLH+we+xw/rNTF8PKoQgEaCD4+hh6WSDlvgKyNWFvrLswXtGU4pOWlEex1pweYILdFBH
ypKTFFZ/2jmZFTgfnjAH3BWwmx7p5kcrmESVUgnkyriRginX3cJqeEXpQuKLdTmJZXyOIDdbpeGd
cg7ZE09iFjA8nq30NbLkJ7SAWghFmxUb63vr3FLCbeo05f0B3F/m6jNDUblSL+BBBf6xlBRqHHE6
EkDZcTYenbteXV12fhFg5a6y3s7a6Rz+ms0sFmxkKvJP2nGu53eRuRQXxkyd3rKzXJJEupoEeN+D
HznjHEIqYxmgGYoST36om+Sf29d8aU03ZHjyGG0q0/3MRNbc3wSEYD4rU/2f5wEIhPi+huXuvy0x
0Bgyt7i82KzCmV0nflWXSfaOTK2Rgx/NYXmpQqAa34xLlQlfuAz2QX4r7uaRtH17lvd3y0Ugu5yz
gdp3YYjipTR5bpvXFsGuIehDGndp45tefyTmMPl/K/FPc9EoPdL7Sz9DtimQQJuGAy0yd4YJixSd
CoEdcya+eyHTdqu6on0XYan3m2+ggfMrXfPXmJcamlETRXpUfiXL/WBEDWxoUH9vckmZ2sXnE3PL
BH4J5E/JT2EbR9vN+qa+hSAy0u5s9lYHTng+l8Y1IWnOdAdVPl4kNylbiEQYyTj400WCo8lYzL7w
rLYghMl/NYYwvLuFWEaqjkL3l9n+TdF0AAz3Iwr23Gjsy8/X5+h5RygQhYrfrZgX8Tv2thhbX8dL
UqVBxSWuyB1R99etRwxPAa1/roCvviqbRyx9CO3abAnjvQ683jZLl+PpGx3Lo08JsEjFIq6ulyPr
jSO3Vv9us2oQIv4Z+fbAwDFkDGf3GrK480rgzMiPWPCRxTccjNEpcakCFJbq0Om/lf1OzrM1OEJT
FrykWeSO1L8/cSb4CQ6IYIWzjn3GxbuKJUbneYIH+Kn0t9zxyg9fIKwCcDTWb6e4AVxs58lbKpRy
zGU00H27k1v61/gRf/XMUo7x+dlYRwH8UIiPjr5z4XznRa+Mt9dDi7orqHo+msEa/8qNdw0/DGYi
KrkPf+uw7HZnPlnsKaq2apLMOqrV7SHSkPqKtfvWWksdW9PL+Brq3bzP8JbgXKZ3dlouyz1kiZQO
5kAGUreMvOtjb3UE8G4yNrpVEtsM7IQresfs6pq2M6HuiN8Nj3O8paEsTy77X0l0Jwc2UkI/GYnW
YszBKZVlBcapAdf6tfpEvirZrn9dVG+K43AcQQW9BLk2dXK6tN2nTxSFEyKnFTjyqRfmrvvgVuyT
uEJXPLJUo1FogLw5+aomo6M92QfpcZsu5cITtNPcYpKAC/19biwH2BWwk7ByBeEf2Jbor5zYVvQ4
nma3ojXUtF9XikU5JDQlzAX6NU0GD5KyCk6/+p+Wi/tkDCSVALoxexrAXLeIAHccKsIf6h8f22yW
+i8VU3gFn3bCyKcIK6opqXzTFgbKQ2rheWrOH+Y2V/eqObf1S94w1aAImhC7gYEYhHO7ev4i+N79
l71UXZCzwdp/u199Tms5hp8DAOSfTinWCZPxcXLOpzx3vvSTy3pKO8PfAkcrDz9MddiGD3Ted8ic
DbpDD3xpIWwKaY821LrTmanS3ct1c2CaBdeCWDqTd2z0funMP/T4cbpi4TfSFGX9qHv/XtRuv2qI
ZM05YWQYXSY0fT5cbX2yx8cXNEmhbEyN3dwfRK7zwGk1G0u7b4Mz3TwDHJeNVB8e88Da6VUyopxa
8Xmo3PBnM4dLHyRqPGKXnIBG3PmJtuGmmP5NUko5BCulXqrznP1tkqriCQmdwQOB2QXc2exuE7x6
6Q3mBrv01iEyHUHvVZgF5M4UtGe+LIqNeh39DKMsxI8H8INmYR1XA5mLbsIh6AJBBLOgiLMRZw3x
5fYtbb7ON/0jUJT0d28BUxLsNa6wjXS69ltGbH3pxxkJtGXOYpDBj1TAcViBfLRcCTlZGB7uDj4a
6scYPs/HUBWSPJZlqfi81erLksD2NSOWr6fLbT8XofnvzC16oa9rjecXU4duH98nYbxoNRV9WXcc
kHgpLDnP6+YGVf2Zixg8oX1KjqLRoB8J+idJFopXIDjyOfJLsLbs0+KAfI51JmAisP/T4ickG2zA
pVlZ/ft5LMsWVsP3aC+pGf3RFcWaJdIHktyDXBrvz5MdOLSd8xzW6h0OtlpphjcHqjdHpxuPXZVE
vvjzOdPraguewbRAhiMn3mvD8tL9zVTnGy2L7rwcwkUVJFOeRBb1OyUDoafZRF2zyTmghmTSYgyU
hxHrZPZX90hdvW5d4spkTs49K/Tk0Ol8mt5vK3I7as9wRbx0Fsol5WvyEfmo2VYn/WSBaIyzvCdO
4uJFyjNiEvrCLncHWB6cnFmEtxF9Gk2DJb8sdEBqvprd8xYpmhVlnrDpxz6P/IFKPnbqOPPuLxFh
DF5O8/MmIpytVWvfsShXDUYR5ZxtYpSZTLc1DUiN9+ZaMNxaaXbFUdHDoOEhFLclb0M85PB7U+zh
EgOkd0j3o+J/y8ODeDdQ8e9Tt6OMGLW65AuByWn+FNopM0/mIxSLtF6tqfr7riegxoyRJvDiswy9
hE5h+M6jMWL3jaXFtC1srTiAnRJzoxIxDHthV7ah/zkHFxSXj5bHuC/Wi+P04MNiy3YcPpTvHjfZ
9NjeyyFKNbT9+N1Wj4TxeMd7EJu/U3nvMCKFg6lAyWPdCgNoqo9TCjRdWKKpUowhRaHvsWf/8JdV
qXcugyubvAOLOr4iy8UndX7zQuBD6k8vu2Ya9gTcyG/UrkvOFxOIKDXlXhx3/GGpyXFOIW9kJesT
h15J3KwgWJ6vNPPlw0DwcEChbKHNm+HmkIu+3Vxh3uH4N+ub6wwwhcEH5RPDc9Xnu7V0ujUO4Ufx
v+iWKhbiHJpQBwvQXnuEaHOa4jhq38qLwdjANbXctcUH4SQGcKhZadmJ7EDY2Zd867iPIrnmTzlF
4U+QnVteasiQCX8+r74NWp4ywHRAanX8jVEaU47EVGSccwTzM0gi+a7C7sXwgRBys4OIQahejzGC
vb+UaTsqU/pS9KMkLjOWmICrIrtIvhFyG1qiMGqm7nXEEtmJB9aZPmZPCORJ8jNWdtF6ufQPX457
Bbu3Wih+kzBUk6Fbok1tPcDXlZCHCrRkgbWKt0aChpAp/kvYYicKd9lTKBfBhS9U8H8ld5YqiEnF
99rvppZPNhmUevBBzWPAbN/uy4vQqoX6AY1IGhk34OO6FcQzq+8IYg9cmr8GtDni0o0iTljIpNl4
h9rUzkZH3/4rYElBlEGt2vqmMhlt5bF0Ryxlc1NxbE6jl5VRnlVqe0t8xbpd43n24NogfYZgZ2x/
mvFqNt+8kYwt29zqEEaLPKb31YQnKfFoSjCd+i4UKbx2Datzq5PovlMGsbYyOKfWsfYAxgJ6LpcA
hXYQHPtwAhuKS+z+KJ+tKvneAGNc+xa0DFS3ACG/VhRRn/q9WSWEOVrh+XX8JqhwLgfX/pqCPVyg
twUpX+4lswTWlsgP43RwBGGVh6OD8OCWEaqS+bfhylKgHTMa+jXRx0tGSgzVWWFTwuI7BfNdpvQX
A2XqJqxVWPMg0+LUpXlBalAXm8Y5lmusgfpEIx1Y9EoKu6tnC8EXWNfHE/ntq5xgPkpVn6As09+y
dJL7ITYi22twOGKfsOMQKYxwVmQdiR9eEZk2rzb7Ut2dHP4vojAVkxhCv7nxSxmhaLAUEIWDi4LF
uDU7VVhIiUZgi8V7OoSG8LhCuvFO5y30u7tr+8UpHWQrmgAIleIU+yBDGnzByZl4Xf2XYeW2S5ru
qvf3FqHnP5hpLldxiks5YMrdIcd4fVFtfJHQPjJIFnv/a7L+GLeGVYUMRJHoF4AR0ptzY/ze0QYn
dY40aoK7m14guvCG9gTbOEp3CsJzdAsXgkLMOvrmnbbAjzjAiGZXNLzMk+zUZ5hNe6+GK0CryznC
ArjFOM4y/tvqhxhiaKsN+AS/tOjhY1i/E/WrYKy4Z2hYM5+0rUXO8i48BwruzESPYko/3jWXpGNu
rfa6qQr1DLzpl1V7NFnDBexHk6xdZ8eh3Px3L3D4EBFac64POOT9+VmzDinhrWoPHp/ePcc/l/l5
G5G/VN3cS03m6G9rVcfGkBbKl3Kp6dgVuZmH6iwh84A3KJgd1bsk52TYf3H7cRXzbAYnlGRnPlI/
m/6c+W8JHuu2q/JZRcy+2OA1dU7nNj7+dUl2FyKsy+J04LxCtuVYKD7lKvAPsab8dPRJ224Zrid0
xkyvNWu/eF6hCg/D5GqWBSjXwFOyVAO29eMgn5fSDOX+iLOt+lsDeJsQCS0jBPx8rLs5QEhihDOb
M/bxEyxYjTvtvR3wMysrnIh1HIsf1EOsw9eQgoPRVLqZIJiXkm7yrAtGkA0ec5zFzblXRQV/0Vld
mPz0S219x4zGQKemkYqAHfqCgKUKasyN9kQ9VyEe+xhnZDxgVBhtUqLonRor+TOX8x50aUOPYzAS
CnSlT4iGVAcgSU3k5Sn/DzFYTIrJryDztqcpIA5xV5T+GCItktM0JiMLKM4xX/G3DsSpq3joEB0y
t22LugYw7a5aL27KS1mQ2b6czWEiaiJ5uz6r0Doc6bZ2DgUx/oeYScsXviRwCHrxGM6EgkXj1cf+
9QGCnXMryn9heqXTCaLkxBlvnai79cy28p8wshIN0+BeiYCLRKr8+UfoD8MLjgiPYr6Gq+GDJezh
6+LkuddJSJhKcw6oLeYHCDPXCJozXjfu0YYsrUfoAehp/hpM9hhAbCpXuZwGaFwCmLdJtT4AtXqT
oUQLIEXlgfJQ63kMWPsawXfFSoiI2lw97OaZdx2fQHxN/eqdEenGpYR0RqSe8qfCDZUqFUsQg60g
llWA9OXPHsyeJ2wOj3hZR+JdioMAU5FBf/I5+XZTIn+eAdC0Orkh9NX8/8Q/tArgB1iOtc0NPTS5
OZIOVgmzgco0kGqA7kloxQsXieAiD5+iesXKfpccXRn411vBKy/h3BhIlO2BCclvm6YeecT+VNX7
GZVKDA9NL64CZwIPQ5X086aeTEi6nMGqkHnADIiq4jT4sMwdS/HNtmGybXIU4hEguUtMobOhwyK6
Nf+mM+7Tj6MfRQZ35v+RUaP7mkhw4z448+CDAuwZsLeTie78jrCTm76fBgn0qemBhBKqXgfD+SBc
6AGaqL2psPeEdNSjUE4bprnNl+njI4MKqstG5idbg2o50rfsMra5t+2SMKrvVU23lD1Sl5icL3Tp
1qQCvq4geAC1tLVSNn2Ta8AHphEy+3EH6TkIgSGK54BR6N+/h2M2Wo4z6qbXO6bcQuhH8doi/jV6
I3dWQ80G+hILoulLkyQatN0oGNHQ3iAql4xPMK44PWcm2/8k/Z4mKIH2ccEkg8lH0Lq0KW8fDtQI
ZcMKI6eTPl/U4nC+GBaH0wNm3cR4mdbRPYW6Ek7/xdGGWsBwu+uOyUKHqOvFnY0DldTS8O3v6RnT
1M42/2fmYPN3OW6/mGTnlo2E4EB8TCGu0XkAY2oBuU+ceniNOfO5TCJ6TdC7HYQFZC4v21U2EDsk
c+EKG+FecSk7rvYzidK2Nlc2gtGQoJT+jSlu2X9pmiz5a1N+VnyoQtAZVPtEczmMbU6YZkCCZ4Y9
S5lKOR4QpPpAdrn+nAwUGRt/KCk8iCMENEHbKnBjD/8wFDoDH7KqAABQ1lOtVs2St4EJBsIYLw2u
YAg1/Su+R++RNmD6+tKYONXEafVOr4JaJ3dgZFGTUOQJSrKiyD9eBUwnF/NUMMFBT0n7GAr4Ez0l
vd4aEvvLQznYL8UW3kKfpThVsmgnx5ySPo9oV1eTq9PC1TeO5w/KacNC1QoBw8eq/hE3KUn+v7ql
WVwHQ4qbFrAHXzn1hcIP+CXwcEigsP27HcpamKGKRa7CEi5jQN396dyDEuq05KUfanPbbmT+o/5w
9syOcCTG2k6U3u2w1AoWvEAiEzIxp5bTHaRX2qN+mJibyVkwa1+p37v+gE0XVMquZ48NioGens5Q
9lm2eYXuec3WqKQc1DMb1oJ3sCnXCGJ5lsh56do/VusQ3DGgi3QckhDs3pxZ2hqAkO00IQUFq4Wi
TE5Uc1owGVRaxh5RKSXvwcgHYp3Fd1LaNMB1TNd2+sGFc6pio3PqHUpuyC2YudQu5/HNUUkLiXhU
c7sh/y8SyU472EoO/eE6m8R2vgldWvw0wfgso0UfnBohubs6H+MHypdQe1kpktimFqItIUiNcK0w
xohrI+8truzHLDjT8ifnqj2Qf8d9n0jyutORiRw3U+4Va59XhxYFzjBs4Jz+9GWrSYs0RGW/WLDv
6bqb89AM4X2mj+NT/H7PG3SGCbm643mvrWyppZVolLYfZMGSHn/vzfGNbK/h8QokxhwB785KUglB
2TlOkAYMYxWJ4SdEWeIkrZgX2FGKrsRIxVg8iQeIMG+hbQMB2KSXd6j5+TIGau4liZdVpS6GB42D
Yuc1KdP6W9eX5Xt7BhhhNvpRPMWXJ8oXc1q4qMrFko9GcPggHC4cqHi8wjbP3P0ZNBppOQm2juGG
fZLLYOR0MHY9dynm5l66J6a4jwEy7us24w7ydSbKAXUdWjMqSUWSKcwdHw+GVaDMaAm0RS29h0YJ
pnSu4PgJn8SazWljXQjQV90dZ/xx/mEg+Aw0FxPMjdr74tkq7bfM0E2bmNSByz9O9SsW5XzhWFrX
GcMoT9l49tO6iSp/6mygNdu2oVLTQbw6H+0zQ7je5jFo/CG2Drad+f7voreFurASqQIGuhRf8h4h
CQCwI2rHP5vr0mE1ja76ZHOLehG8fLQvF2S1WCYminGedrIzbpPUPRmaszi7TIVoXXhVQ7mmLsaq
TNbqxzwfVXGfuCUqDI3oK5NtSVxEiCUAj2Z6Xhh3xznAocIA58NlQbXHxVRsxg5EnNGNEeXglKB6
dAXnPQYOuBKP9JF7nz7Ezaw7mbh8LPl/OnvsK4UbtAN8u7nIStlxDuOYYKpBf5nmOFmfopErUTLE
SPx9xlEj3EQn9IU1hHDijtPVWM/ej6gC1hU77VLfw5OYOniushKP9OJEuJ21pIwpR4c1SUvExOkn
2ji2IWw3sPo00siO0BeQ8YNzGIPPblbZBzLxIXR+ksA+94Rgs6znUB9C48wj95HJEtBl0pG9BzUy
xoby9TaX7jZj/DE8Eu18+FoLDGYw95RIMKsr9XbZj3lZ9KxN89gLgD10gxxHYdzPQmI9pzf7YUJf
UyOALPMWAEFMa8eZNGKK+TvlomRRYfuy6zyk3pU3wGUz4nGcr55tBYrJ/3YKbjSiQi4Uk2P35Qw9
M975pq/Y6oMAiW2WpxujHl5h2KVDwTg3olzh36/XloV1W8NYY0zIRBpfEBAho4UZ62ATI/3SZLOZ
qiYRMg3HeJm9i5EdfKwqQntM0XSh4wiTIf+xe5HefTpohKfptJ8BXnPZPVPIPl/BzK9JJpDKV4lg
I4s6MPyuUozKZ0Y0fUuWi4bflq035UmY5NzLItLW697kFa/kRifzGQeWTUkjOKUfrZR9WoOu2iYy
tFxI7brjeNWG/Hdz9D+EkHrU4GZQIK51BkjXycg84c0okpcLePLi8HhOTROmC/6fYuLuinm8msd6
eYxv7SaKoaTEIXaHaYyzQBqqzOoyL+hqQZs3LC54NHaKPo0g3z0dsUxzNgqpZ6kHnN7zf9KttgD4
WZJMKeorGB4gz44qDNa/7Eypyic1dCfeRnJtBjsAPvNa1FdhQVXUJeL9ZhkrhSyv2qv/RJXnWCPG
4VxA7PJN1kwxdyh87Od3hOTe3AOopBBkFNwuZ6bHavzDEQG2tCcyqY0kfOWvp7fEbSBRQdlQINd8
D3w72rKW0y1txFAAgkPqrkn82tzkE0P6q1rbOrL9IVQF2kaQfKmQneUTo/tFfy9xJTRoJQG+Ikq7
VCQGrSaLJ6EChol/eXJoqRuDDLfNBm5aXBXKfeepxwuxN5Q2IyLz5VsEz8E7T2HbqXVbwAgnPMB3
oAGcL0oF5Q0B92OTlo+Z3SxZSAyStxh6jJ2ur3wAbfGz8/P+ljTV15SO/jYCxxAed2aHiqUjdCNR
ozM1tLJxFT+jHsfW0D8OE2oLIbaQKm4oc90X9Wo1B5UcQrRRYaOCJNCsGBDT/cgUjpVO1/kwFoYH
T09QdDkC+7cwYSFV8qCorBr+0KMvDNaTLpJG/gFcboaHh7FpgytOkiu1wMtDg2Lu8L1EEAiA8Txy
XP1G3D0s70lBOcD4pWxBIyrpBrNyJlMzEQ/M0eb6Xa9JzE434chbklWnzX4pj/OVdrlFX8JKFfYE
1PH/keryCWBRqPc5D6HWaOWwl8E8PxzaGtwtfglU2NPCvfZ+yNY6ODAU9U9ZD+MOu1Ml2x8znqi2
E/hl+vXmRaBZvKQNHdF13MnY730Cj5wrleojlsROON5LaS39fIYjL/ZqGBFOYw8c1vynRJNwDDaP
0dfzfxt3T81ui4FqMKN8WlrYBOKNjjwf5bfNDdJS9mZJdIDJB3gFou97bxqijCibYjAMR3Nc7dRs
MqokSCXFrR4VEXd/EY7G5iaJIXFQtAtzXK1DYNlPo6e/q2B3JkUJlHhUW5mVlKinNVbRWCE2lVp+
akiIMgSV+en0ldsc3YSsxp+Y0ghM+2q9BO9DwYIMbd1iP6kfpMZRh4h7syfea/T7XdEjxJ252XAG
p2eZSEbEJzQ+R1C9OlT29nP2np9ORJS/NMRED2Nz8vOG2BVbE2jDZTc4fEp0ZVPCQPbBxbFakamp
xQp5kofcepGEY2y5EiktoXMxx+iKJecuIEH/H9hsZq2wxhtj6C4b8Rc9ozOrMeMAvMukg41yO2Kc
HP+UheVMaEhU2YtIFzfYOOXFOYPJle0MpaCinF98da/T16kfWu5UAnqbiVtpJJ5zr+ufqiKEbAW7
IDuRQiINRqnPgpbHt8Xlr9sGzwAtYiGemCMe34EiuXYEhXeNv0L67ELe4C/zusXTCUkOWQlxwtry
C+9u+pxT8KyD72Fan5pWUqM8OGYx4x31ZzigUN0ntL2EyzgVnBMmOISgiPhrgl18fp2GwZ3j1mxL
5XuNpfR6lPeS25sh7OB2t6C1bVw6a5UFq1CvIcMjbC0mH9bykIns1QxJ6jRicLJr15thWUUhe6oe
iMGqd8bprbTURTOon/jzQOryl71tOnMsRJ/TxEpffbAX+Zfx+qO8AkFUj+dTxDDoC4pxvuT6ybEB
1XJ2TMUSBiKVb7gcxFI3rsC6TaO+i8FvYW1jSneT0ynlwTNZnUjXFf7hk/+6j8P3Oy9JWA95H52H
8wQnvfL7KzcTsYRSuTB4A9Qv0iofo5F5RlhadQVkaKoG770iOqG1csXshZ67X2L6XzjK3uoWSYhW
hSIVTKGGqZjxhG6S3b3GJ+xziwUbkw9LgY6tedDPtuUHOcS/7CgSz07n97DLANsCYdtwuCgHZbWc
BKT06CKJEio8vqu5z9jqKx2PVJfLWqQy2ZpgJQZu9ZNqe/AQOKlv6pYDD5Dj5yLZvvEClSsFysIq
4Q34lPKXu3u+JjMyEJ3TFoOxyNlh4pgx2Xi8+JQYSytE9YxFx4upE7JUTehbhJlkz+oxyP30RJt9
0RxnNZOkiCH7t5DB4LSRwraIrEdXVYKPVKR3Qxr5h2aw1M3jhUQqFFRvCMKb4huRsHhYttdTSTJ5
5KiJsmExF135s0d0DFr7mS6sof3O1NlwtQHXb+biog+Lp4ufSidUUJ/jn7Uzkg3HBbhWu7x2xz9b
rWh4Af9FQOPtujCIBSVTPaAiaHATwOxd1nDIbrGgWQnARZLxy2rv0pGTUzwPLedv7ozYxTmLij8i
y7D5tmWRDC/2KkVlTry8qw9s6lM0gYiqEx08bJiW6SLHqnuI6BjBx9+c369IUM/F0PFSGzvsLHLv
MmezC6hokOYT45pIaiXjGSTzuala3tf+j/B1Yx/QvlAz4l0ljyED25gAyb43HOgcOV0D7R2S0x4c
mbOvcE4IS2ZxyxeznD+S2tZD7CyjF75ox4DZlmzd/6Cvdj/wp7bJFMJI7WZiRytv0M/+bxtTQ1J8
J7BOVH2ceXCiSuf8fvnUZFs4/D71yRt3ct0GcvyeTVNH4g1lAON9dqW8XVuth3OqFpuDaeLGpJ14
CtZgBkgOlEHjZyTpOQuLXgKGRlbsa3h1AuVItAHrB5KwvAAccj0eIG8LRKqFf4acmeBNl42eGtzs
aO8/corIrEeLF/fOqQCYdZY+2HqQZyLT82KxTainpGIeH+iIrp3mym1flJWWYsLJl7vjwuLaq2sI
TG2J7L2tnrzxoIRhhjclMF8M81xMmBNJBm5EWAkifZmhQqnEpD45AbHz7slJUsdCPCi+udOhxdUi
PbtdCAtLIvkhGIUgR9Z9VTDWvoUfvsBHsBvgA1hwULNOCQEn1csGwJIbGRgBOBrdmIN1OaSR9WDb
1yikLpeK16DeA5JVAQVOOEvbZHr/ROvE86Gbb5Dbae1zXIbfGaPluHG2pLzUd5Sqt45dcPQ3Ys5/
wXVbadR5S+ZSCM1g2L6tgIj36/BmwG9GZjvnWEXbR5YMEiVS+DC80gRrpRbFuYo+iFQlicajwbDD
L4EUftg4EKKkwRkNZjIjn+M5SEsymvGN5Q7/cl4dw9dus5UVt6NP518F443UvljWve1p8zE2gkUA
IdUyDzJwczqakTnQppJZLb3hJSQlbzlCWecQfxhS6QnXYd3jYpEVHpvlZe5nYrAYcM+pFSxBTlYB
DubytZkanP4DuI/LI8wVZVqywt/HnJ8+7f+QMdStJVXHrnQQyly0isGhntAxl2M0PuE16iM3Ozm3
hT2QM7BJQ0EKFSYZD7BWH+7v02xKxl3mR6SfMhbO8U4/8NwHlfycs4q3I7MP9lyHrD0b/tyyvnCV
FYbSdU1ul4iPwLuOoXb4QtsCIlSEft9KSxho03Z5DJVoNJ7t3HoseVWGSYFe4n38j5nRN5i8RtD+
ynezGeUGyPgGKr7A9/xsHdpMkZRLFm/VL+93DAs79gMIhlZxG/yDHX/JRjCJZFbIkDF9TITnzzOC
QowXyRoPNN678LpQ0NT2OI5NocCkU+GvrzewCKYrKqsHohF3aaCq0ik4HQZPAe1uDPggJ+M1ENMs
IzmNW7xadvMmaDb56Tw8yHltiJDJsBiE5V9v+0IkjY3IHONfN0WxfjSWs/smBzkAIIP1LMKMFyXo
1gLQ7EJqQxsQMa4WqsIUjUQdSiKhj/coJoxGQFsjQc+CrTZZrgHCy6ohGK8HVsfk4ctNQezcS0LF
9UZeIjnA8+Xum1v68J90Q9RlpKyXBSWUNKlJHqSRboC7G4OMzfCs4Jdth1YNZHprrFVtBjE9wmTQ
i0o4y6kPN35Uhmfvrw7ACKBBiUnDu/n9D9oXHeULDMTItul1BCguRI/zYwrhl833Ld9+HhdpHbLP
pACRcYvr5fsI3PhtmhlUWjTK7mYtCQofic90K5FX1DpdLOPduqc30nnRnD8RN/mmShlDggc/avef
m6mUdbneVxJju5rQFMQ7aWa6ga6YI2dWMBO83bBRlzPDiyOsDSxilJHfFac6+XPVE0YUknGjvsMg
geBwUgJNrE/6o6PF8xXMY0+bOWQP+1ej0P7XH2eBd0+AxtofeKU6jzARe4OpL7xDEfDJiTce4Y+W
gsBUnOUeZD+njvdORGaj1r1hYFVliyZO7VNmQ7t06+NUF2kWDr7TmXwrq76ZrKHZCz9y1cQ0S+x7
eydw1rauOzBLWlGn+Clw3jWvKKxytgXBw3C2YyZEyVbA9iREML8WvLGys6zrSXkQ6LTuZw0ImuSB
iewiXCntCRI/9pXHJslivVKLg0UkbCs5tnCsizIIfo6SEeY+ppg8IDQcXVC4Ay+cYE20cf9R5qWp
+oyizL9kRAK7wzN8JYbdEvRrBZ+J1ZB3l8xKHP++xRUhu2wAJDYkuPntCxB0E4r6IJycl/oSpa7a
D5y+qHb1jAaMS5UlY0XUaahPMc27VPL0PYuVdhGLYhX34LDZpkZVSq4POKCvc6QjM3aaLOlLCl8s
HENG8t2egSVowjM3/XfCJ4YQS9u9xEwyse9P2p++bhNfyNEbhoEFsu/CbScQGeSsZreytQWShiF3
R1x8h8EKQokXUfBfxSXw53vxIk51X4XigEgJdEcFVyoWuPhz9JEavX/fIrkNp0xbUNqQJ8pS/7sG
YrUbsNa77HQH7kolrbOE63HnoxLhsj0fBK1ToawOTcTIqKFsAFyhpZziZ8aLc6y28Fah2YlDdmPH
VS4IPj/+rJ7MtlLeDc11HOmtEx2V2CtwubKsJtiY+kAXi3ieWWTF/q9/9qRxJmvgTYEAUoIy3097
8Z9+fmzVxTThaBMT56wLWpvPB5qvJC5u7hbKfYo6PPMgWBi+GyQ86NgBrT0eCFrs/cbcF1lbAgLK
fz9mbdeQ4bpxsPdLDrYPVLDjwuLFJA+JCoNQQ2cW6napig2l5FEd1brJaJ295JkExZgLbkxRLBoR
yu6JYFUzhH0sRnYMxOcLbmSNJMB5XHSEw9/TAH2tXILGjjTWd4q1S30hpy+9CFlZwj/SonZS83ib
iRWbfNUj9U6sD/HKmP7asDbIfnUwDcCISLvepuZe6xwo2YbIBjGsHDOcUNy5EB9Axkt8liR5Qef+
snXTW9OpAPe93PlYbvR5u7yhKQWnIhxQV7iuaSX02F+F9mXPq8P3vtMSxiIpLQVVM6xvGIT9zcFf
vidiV/jbVoPeIZrIZShM9EYcaupo5GjQ87HeA0/QPbY5hitRA/Qtkrw/pfJJozH7UyINJtYSdHr+
HQLLrWeb2gVkvQQJ+9piP9RAuIycCc779AeCFWpFcLklK6suojVoPeX72INJvrCPQdoOqkldp1lH
ii/baYz70Lc7IDnkVgy2dnBDmHrr3uxX4XGzZd9Gvk3zDHn8sS9dA8ek9A6uYEeOkeZd/CiP+XOH
ECHR8GpoirMbDxBAfbdEnmfMKYg8G2SePLX+l3dcTTKvlCwG3/A3fyJUV9zanQZXptQnneGOn/Ey
a8a91sdsM0dn2hb8G9AJ4rMzIdcxo5m73TM9eXKYD41AWuge8IbDFmWHqHrr5nJCtbNLUG0GEuOg
n6IrQBlS85AiU2jocQy5HQJ/OzeRlnooDH2CkcZI8h6oYOzd69y24cK5MNi4RFaDdHx/misVn66X
I+6ie0vd1u0KwO4ha2vIxJ28r4bgjywMlMTXdCPXCxh+lmlPRuNQbWjLI9DVKmodWJR9pKSrXrnQ
aqD1O71MDhz0Bttu8KyKXcWf+Z/87LukUfBti//+g+ejIEN7fyBdfpkrsnzybYsKK5sFIaBxGAIf
sRdVhirYotg+Jc3s51bEsHEbNv5HsMiCG4I5APdX6kqX4RI7E383QK8u6etxqUyrj+xsvCPMAxri
MxZ5tCNDadPnl03wjGWSZa4rI7dKG2HnQHwTi+RfwGBFx304qdeQ6TU5BPTyokNBn4Jo4zAkN+4I
+ShuADiA3e0hTIajC/QwaodxW55e6vZQxXQgkLADSYrCRHBmwH9zOFCcy0BYBjoLzLH6lsVQx+Mp
7bjV20kiWjHWxlcttBof1Ddf/v+2wmAX1bZuBAC8ncomaVazCjYBrUbXXSwJrCYEmi3qIDbWq5vY
poCpYM7fJKkiVPDFA2sYTU4DB47sggda095A7dLaaeUQaXDpJp58pavQOy511giR/frVNyyp75+m
CaYU125K+Ysle0aiy4bEiEjnfN2ZiisofXywPN6IK+NQ6K1jy2tyR+ChVTJ3R+F/5uKFKMQ7Jev1
prHeOq6bx7fhKGZ+0TPGvY/HxgOGVpCegrwuSg6xoPRwftiswAWPHRxw994GDJ1hGHNlir0uX5Qa
h8xNTbKBhJqaKZ9qgjF1sKpywcASkfu5NkDf41tZpkaAgKtHQENngKsvf78oPUI9avSA9QXpTG5X
kQe2Kx4QZCgkVFwKSuxJtqVKUmPtDSj8ywi7ZyENzcm/GSWdu7VPZC7Ien5Na0beatvYNZpY2tup
xmnVWON2joLZ1GSqFodQC4AzzjEnUyr8WgmP//W4d8YsZIKHLHTsOLmCx2HMrCkySY/0EiZzgetc
aA0tBTyfviJKLul0tKMeZfrkAB3RjsMCg20SySnT5g40VHFBMg8L/9ypDUSh7gDmImlF+zjVjGx6
88njN9d7i1EBgMer9+QAihgrWtSQonbL278IEpIjvGjLaxDVg9tjik/w2zmolDNVv2RS34vBHcrf
sDqzAkWSGe2UgZ7wzhlC5P3dwO8BH2k1TnkUxbz6qePY0Xxa4N+PTlXEgbeokwriZEHePK6ViDTx
HsCLftNChre+MnbkDF01q9DjuGQy9S/N97AMl53z6FnUOPEmCcPNhPog7ZbOmGjEkgkbLSKu2YjP
TEWFtnU8lODxGCimg0RgoFzClnzIFqd7J477w8ebw7ts+Ww7ovr2q63Mg/Pa8Ocu5OkNK3jAb790
eSc4dWI8Q2ADqUhcBUdNtx5Fwr22Lu/XXePMnN7bxmIhCaCmmrCC6DwUXafzWlnqLdhR7ooPOvya
UetGKw0q9He4f3cXuajGldJVEE1oET8DqBf/HSvvTaXxfqDsk88YiS4j2xZw/GLsfmcX7ow1Sc9S
ODcS/U426EsAI5mR9Fc6ik3cj0hV7/l0uh6P5l1oyfMSN0sSPCABeK9vtNdmMYt4Sa14J4pjFLTL
dyc8/iGCyfN3gy8e6zgmm9VDaG0okxKk5jFbUctQfO+ynEyrFPbJpTMaZVI+xjlKUrb7S2CPVggr
X2P96DdCxDs/UE5EC13emHMAQSl5ISrECNEAVKk8BV4SZWZL7CgYUdAQpza6sLgroS4HCZO5LO4x
k+DyAK6DvsBnUd5b66pqYIy4PDk+cK3FObCuWyg+qjxE0Ccr9J7orvlfhJ/IAH5kmXOJTmc7tfdN
fle3uz3uk1HsWHtSh9IRkMPi6lktwrsQOmn4+By9+L7ZW4LUxOfqP/y1pQGL+8mXNSyPSLS0i0IK
L7jMXKoC3udjacGYgG6qhOc2dGdjHt4gtmdH0FHVlTOcyNuVNrtKUDglYECnK3V4j2Z83JsM/+YI
tHLs5mbC3ANS+WPdZlDfJAlHbjkUpdXOG/VL/ipzHVKrCvH4vmyrsGgVsPXcO14AQsJ+4R48xqln
uvdyQ7KpwC5k10RVLoTLxGWvfxR+cyqS46o2GuVPsdHDWse0qX/G6bIMn22oggHD6YIpC8ZvLWUL
gKuVVQyGAOSJWgsUgZdwZZDcdcKQWOc1M7rPOC85ynmX/G1cG2HgopYHwu7ZHw23XEgJWALn79+6
I/4719fY5EK2Z3N48Dkk2GYIITa3e9hSxHyWGWUDX7J6hEHJd5/OUQDnNqryZLFaL9RJG7kEJ1jM
+PwAl2nPXNaLMKMtoQ6NR5sVkm6qA6tZc5e3bWIKvJ0kcxhp1+s93GtiqL8WzCWoYXIJxzLPVNqk
prbH8lZePXjuP7m5OBchGMeb8ISMXyASN38hb+snSYa5ue+7WH9ttfD+lEqC85YRAypLIiKUBOj3
CTNEpe6kp8gZ0V7jNzSPng/VPx1ilqE8KZgwUzElN20kYMFdUApaXpgTKLxd2UGNNJjFFd/VdXXy
ZZBbKmfbhxspH6Hi01hVVO4dct35P8gJtRVj68I4Qwf1JbbqT1g0vgh1zPH/6hedS1KUkpPBSdg8
ENxkh8QgrvxtuXDV3Spr8mB7xbMt3Qg8n9x171Ueq25u4a2T0ErPnxz4xKnqywkCqjyL4Gz/YCE6
IxSkh6FUC87jn0LEOgvlHqDTRrcwLn2g32MeRvCChEyFBnXk9vKThkp6lGrMgXwAU+ukIbRWAByd
ctgnnrxjIevMoZzR2CyDepBnYrtGEfiiUzbx8VOiEIj0Nbxj4zSmJ6zBSy0DHYe8+cnL6h83lMZ5
KPs9mRr0rr3wao4f3SDMznhLdFp7s5pfAEEReZCzu8qKMESYkL7TPl+Rzo2OS1w0ZL6HXbjAqQjP
U1Q3WkHM2/hZbELoyd7zqrUEtDbx/BAZiX1KI0INRrwHRAOjp4r3LjSSR2zkJCqGxATNM3olxF9n
13dxDLeUy7EWVFWRLdlGRb68js6P4VxKyM0BvVCDg4qSNsZCgzhVxSjCgf5KMmdksUHKGLPWjyEk
GBrbD2oTNRJzDgTvHsHy1W0anO1yk/I36RYzz0mHvOWgpUrfOybmtPRdDzcMs4ohIioHr9TkMNv+
2Tv7KgCGLV2rJPartb0GfPAQ6XgPtrz2JyG0f7saD7LKd6Ps59sHbX0ct0ws7ANFS4Ax9cdX4KYi
CiMwGJDdqDQQEUYFX9P+7b2Xg3DoZfoBqWMX2YlfB7gaDzQiWqUvFAja7j4fksZKTS/jsg0XmQXV
ue3Dkpuo7hl+v98eg9/54Xv1t/ByNKxqB2iRZI6a54ROyPqyRZztZ+Nm1NMXbkkvkicXMvoD09Uk
CUMbyv13ONAgiRXUQpVb9sCLWifg5U/KhDb1PcCNmsdmitupLDNIZAUKuBUQ9a+X5E3w3DJViG4s
Bto4txog13mgvORCGjSjSwp1Gw4h3LFBXDzgHBedpmV+GomvfYnR/u8ZBN0/9hqYVe/y5PKEAVfL
9J19YI4IJ7FfPsvhPH3S9pMT1wgI0Z0C+mOh8JxWMJMI/z6+w2ZSwS+/Ovcb/5zJ1JaddnzVsT4r
qMYRlQmopaAYfxQ7u+EZMUJFd80vuFeI+qduIx/MB8FH8lfEAgypEGFdyTVeOSEpSJ2xBrxTnQVc
D9OBwO8YvPxExYe91XyniO6Jgs6154cPaZDOPpjgOVD+nysFtIVLgDxWNCahZBCBaDcF3nts0Hgs
lzITuiqkAVPBh1GIWQU0H9AVV5s3OZHao1MZWEqLp/Hrq8KAkzbdxIju9xOOmTgyK6qD8464ZqlC
Uv5x+st/esUeXseIADuQi9XUbE21mQ5usW8M7sONojhtY4sCqzxip21p2NGGV8xVC1rWl0WvPyXW
jFMpZbPY6W1WsZM9W70CRvLuc9cb43xeMCpZnNQUe3QHpqojaTsbBKTOLXZPSMKzGzq/JNIW0AyQ
N8micff11kMrmyl14V4bsKLD62Z5I+zrlAE/gg7bHXMSLrCDa4hwLt44CXTBDnpEj+FC8FVIPP90
Qz09+GF9uFPtbdMkhbZLkMsIExweXMwlTRno+mXJj6MlKxCS/Y0+Z+3FYtLtcr+vCtE+zUKN0jWq
W1d45eBqwLmGu3QqLEhHfxkpn4q25Oac5CYx08Cq5R1xN0ILYxCvbKEaUqtEC6c4Bcq4CMSH7Ota
Iyh60Ek6NVxUZxiHBl+3HpiJJKuh5GqMtYgmcElhqkEu+P4Z0ksfuocI1dFJ/vDPqDWLe6O7AV7r
iNJ0MvacmjAhxmuF+N0st6xHmCuwecZrXz/T4yDJJByYYdiW0BxTPyfWUlp94KIU3IDL73GbXm5Z
Lyf279gDx17N2O4AQ3P6Rdig9veWdr/O8jRiS/n8OASc/LwxAYuMckBRaATYw21D8IlH4YrbjLNB
cO+nJRHjSjrnxh8L5ZR52HbW7vFNb+fzJS5oewbUSCqDE762zu0Tt2zcuBvaj91CWqaoZ8An34RQ
pGL4M/sdRxfqEE3VFo5+Vu8vY66kQS4iLNW+OSEMincOz/nU5l7TDTfeZyMYmA55vAeVxAlHThnU
JDpUx0yMZfpdp+fPQk8KJIbxU/P0UzkJdeHDIs4UilFr2+s+DojwoFBAXLUTFbqycWdFLjWPzJQ6
Ctcceyj9+L61M89+zhUGDenb5yjv2iIi50KsP/M5yMEJWl4Rs4NUKoOVAoe2uwTTq0YH90nfIdvV
UxmUf7z4Ckm7ruHHjefNC01iKhuJrPgzmqPuyj01tmHuGIZyD08Ed+6zOMcW5Sk6SYq19l9sMe8E
XSK/hIVexSl2IbKLJMC6DqluybHskem+06HVAXQj959h/8PefLisfZ20pDhLI7gEWd52twl/LCwd
2GVtBxBXsLnax8sAofoP5I/0rxs37SiGE7Dp275+57uBrkKJIBcbq/v5F7oGeI7FrxH2XmEHIaJF
3JfQlgU4Foii2pZLTwKe7EQJxyzxVFG83GHfLDy/2yCyzo4jcmYouX1rTGxhxdLXWJ/3CDtKlhSk
0E+kjLkjoBKpQEXXY8ST7UTG4iv/P+xvGuQ7fr+kjkMXXhQIh0hdBy2qB2iBhLDQyHhVKcxd/TNa
0ZrGnJJ+0sB0Hcvx8e1FvysmYJ2u9rPJgCvtjgi5X+N/jLp/ShH9T98B6NmPFUE1wbZeCAHzJYMU
P8HYOkfnvGMjU7jdJ+lEIQ6GcQ2qvQhh3AQzlNaiv8OJKGicnPXAhJbdfSAJ9y35I/BuCciI3XxY
+nmGPpCpbjl3/UEL/HTQz3ExBAwqOAhEkBUkXYhKKM8Yn4LeKp7OADCkFztgMoME1uAmLgS86y5y
W+Ja+6bKJZyS1PXQDIF6wm0WWY5P6ucOJHdWgtwfQ8WHKkeMEyc4I3JgHkqwCM5N9ZS3yG3c/yLL
pRRGanNetk3/J0D/dPbrJYDK4fH/M6qb1MXRNVx1I9O/Nj2tQLe2b/y4D0eH9yYNZjcSFMQcqs2h
l11APlypu2LSUW0mbXUzs4IPsJLZkxy87H/5Kn1TZu8P+heT+FQSS3LHTFr3QP3hTtWnTmQDN2Rq
W0vCV4iqYH3ENmBt5IVpusw3Ge+5DucY4M1Q3OUagc7523a1jGhq/vQVhbOFD9LA6A2Afj+85u45
M9BEnf49xFR7uMeSbw786DzN2w/wfrwz7GAB3VtQfD/fYecssmfRzbir9cPn/x4BHDylMskmd+wS
qrJwuGHjCluZ1Cz66WnPyTTZtNPUIBYqRx4JL/83puLKmH9ZlFOY7f6BKeUbxqAKQjfmdJ1MmJ4A
I4+rFoMPlLfvWrIlrP3x1jMXMmAAxwoY7a/Qp5+A3Wo3S0f41x15vaDvNUXC8tCD8qwU/T4kyMXy
kEo6DYXzGpi2V1sd+GZvV8xdNfbiSAIK7CQF/K89Df7jwk3nQmdeVxWiiz4qVczRvBYomQH8qJF0
PSWqkKuiVTXUrpO6jf9ERPRDAuCJkl5kkea1c/AqW/gP/5RMv57XGRuBKjLvoRSSQwZozTF0voa8
II53T3MG+hgrjxAeUdRAQsDSOClZ0mQJYvmUz2wW2uHLK1JeZHxu4pZHSUfEEXWu/NzB2wQ2J+L0
egXW+jZ+x29MoMPmIA/1VO9vXVB96NzlrexgpIzEvNXr6vrUCCMODpNGrxt/DdbCououiiqXSqGX
Xh5dP21HLEqUNAkatihKqd42c0dG+V9bETcFV1dCiPJpyGUM09Q2Z+9bTblZwPoLjONT3K0+ym1m
FraUZGIXKHg5t2E9fXeUmeQm+xlnJTvfkGhd5u+DyVVhQGUPNuzxjVc6JIVx+ZHbL/4FZKNrQ2aF
iMYxxErIYNnEUr7AvOrXU5PxDtITDzmOGtB/YlZjFQ1iSbp/cAgKREWfRCLW/O5odkxQEWOpH9wc
Z3EXfhUR70cgomkRjAwUqFvRrVLbN5xZklzhpwripOc6JPFOxNN5vaA1Xl7aPALoV6mAoFkSlTMh
et0xJgmW8KDO3dj0eMDuBAT5qQBmzlq2FOmEXc10AmU0p0aOgfmDe8zFEx4EMsQzSXomg3X4ywib
ljr3Bpd6IOIN4E7XE+fcI0Sh09l0gA/vlXf5j7SXTOgoCF2l7HCR63jCth9zK2cSntHn4OQtopGu
Zvn+reHnRoTfTlGAInDUkZRtwB4LzlL/sbOxlmreTsQS/NYPtaE8tPJ3ZZhpiwdiKlIki55hT8er
a8zYtcMlbbM3giswnm7BmYKTf/H7ON/WtzjEcm8JqYo6i0MEdvjstfKApI8cwABv+KtTiWApLR7/
rfTp1Y2Oh6LszbJ5IkwtEnyaOm5YbtK3CgRl6tvI5gT8e5GfDAGXD8+zXU+aMYLlNfCY6+jl4b/J
INy9gh/6i1pVMLX+Uiz3zKQI5rcc3vvH90y9YL61sIWL27i9TQahMNRUdFJlghJop2GotXrSvcqX
EpdjY71Q6PAJ+w/Y7UjHAeCCJb6mrvlGtCLF/c61ZMs8iBJqjo9JT5z5tqi1HH1S/8C0E6nnTWeL
mcKf+CtEcm8fyiHM7VlcJ5elLA9qa62KvmeqrMUYtTnOS3xbLTLm5URZ4+wdYikOG3GXVYlOskip
WE/BKWIpP3FnEgTUmzYv+HEGSJFIzzN9DDkUtghEiml6FSxj3RNHc5syF2D3X0svBDSGgXHTXMAU
Y5Eb/e2iTK75nASc0oZLPohA3sTBUOUVjLopacjUpKBGevC0TY+ftNfvspUQes87Kd17S1w6Q9wV
uJe05w7qSLj/zzcGV0ERFFsR+lHdvX9M75sGIiLderXpfdFIrfIsxK6aVubfZT5sDx7KnPRRsS/k
iVEgMxt9xgwPflRHwPUxWQjqyh9E0EpWMlFg1jvdl7tALX9feCsAM5cEQodB7CoZu459OlYaq0Nz
h5bu7xrJrHqfEJulf4vdKBdfdoeYLwbMAOMffRS3YcaFNHQt0pT/1ZvPAYmPhdoDHyP6NXBkK542
5f+C51nPbc7F0F370xjNl86Uaj749wv2yFbIg5UQIZvd1AJGdf/NmYQ+CCZv0UXBm9UOK+uLAQjG
/dmNugUwYk3zvCuN9E0MScrk2MBNVaK8GTBLYeGVhYcrbhJZ8Y+ipXvFVhe5eStCsPbx6gjvsUQZ
atsNoeLlLVYCR/RPEVT10w42R7mR+A50crjN5taLpQAGvW9h9pLtVJaDGsxXhXF5Tj0WOUsU8ip4
UTtDimeOeUid6hwGWQFU4SKvRNPNLAF7VdCnPdNgp5IWnPpvLHfg03IpZOaRequdHSZIZQWyHzZE
miGduI8w6aq+W9nEN5XLKrHQtaNL+2EiHhKuJsg97LFBNzVVwJy0ilP8DWP8UpdDHBtJP1fAVJN7
lpXQLNZdgbUoozJH+csww+vr2iTdNTvM7Ps4JYwV2Bv9qISqmWXW+nNdNn6aFaobMtCbStndEHvf
rj0j6f0zxultB6/NTWHzfHsjdlQStnq+/TRhDfr5FekRWsDgWF8SwVbcpS6zWhPXxvV+WG//DnRP
PsrATiouJccoS7AFDu7IETbOYbQBo6B3UtHMi14VY3EgrgRvSIZ9jGdEzlFk1F3hVIP4JmGpf0mw
7kEVzRTRg3QjNBSaNaJJ4FVMQIcr5wmWLkyvUXzBM6dhWmAnZEcXLtg2F5P0DwVnPSh5xoycLdI8
hfwfdzB5GLjLfGORaz2BNLu+sTZKfzo8bUsThuLJndXpIweab1c87w+j/LzwusavvmKSN2K0c5Z1
gQF584N++APJgT4WdPOusOjM10dZag0hHkkoDiWMFk0HrAjivhXKpNxxm364QDBmVRuXHkWTPgLA
AcTGQsssH45RHCRDf/6eq2WEHmd2Cmtl1U35ksKWFa4FT6S7iyindKYITyKADkyIis56QnWUv8Ge
DK0HtFB/7OLIuYgXv4IYPpfNaKgALJBYfxd1E9EOcRvVO4lX4ctYn3wLk1A2WdqcE7c7d32U0ucf
VQQnJxr/39q9PKMQG5DFveDA4P+6d/B7NysGGBE1xa3JW6DKcCAkkFsjNXCt7UwExOkj8ktV2mZZ
zKyFP7byIx0cM6figzjgY3VlXu8gpUEz4C6bzLRZ5BcdXncb/JCS7v6FaQOpi5aUkMtbFhVP+WT9
N4JmvvKL/LwlYlktw4096+5RPZqT5zuWpc5IbWz+lq7XqhMkpumXiF7XWUJOzmIxqwDSbEc99szS
6V9a8sz9ViyyDfuXqlwQCTlDEZNXWm0H8YZ+KXp2uLwv7fYpKljsyVMhexefhUlQtV3K2zHFXBmt
+OOFhW3hoPiMzJxGfcz/P4BRIBqSMURyMrSWN5/3pIxD0W/K+mXS+4nUSTeHisrv8K+9tLNDzGYz
FTUmFjdDqx/roTsHcALj/N2FrO1duXSWHAbVzIV/WCZza1wTWhUe40kYfpEioGc0K498r3bvrlEq
Q5wiSRme5E9FkLMNbyPVFJAwbIebWbj433hqKXgJ7uxVzdgtjuPaThMhJV+6ZcJ3DGibL8kdCw1o
ajJQJ42izGMi0AyxWIFCSywKqsNPxoNHVt56cvebQrXoig0hVNcvmQdgD4LSFYCFANa/EOkjEeBz
n/nIVfvC3OQmFciLhBYYpW8CBsiVvzEaQM8hYR+Jvgjt93m10jcMUjimGgRW87/EsUjoleiugE/+
AHbf6ncNs2B3znIRGGF9GBNcsZGh1EXhosKszVDJhcFWlkDMJvIjbCSbHGg59FgoReKqsUcm+Odx
hNYbDAnj4H8c2l6L0wp4PPWHeOhJ7+RwTxfLXT1lejdvnu1fB1q05TOoU+fHVcY+syGyT8BHZWEK
G7uoKKEEqIq3ZgIrWJArEXrJIWHBGaUrnANq1t/14BaPeLrWKc+DYyE52duNs1sbLmJIdK33N/RH
2WhRnjrmBflRmcidlpj/vma72idFv0gmQE/nh+5967PRmOPDsQdL59XjmvIQRMjTHbb2LZjyAEDv
YLgNgBGix/LcnVOD4NMbHO7A8HmJPYlMt2oMR5TQorSBbzExzNwZK9/LOAKCp2+yLV9hryKqfWLS
wH5DyYkQ3TKDv3BTOUJfr5c6vh94seViX0PXhCX8x1p7et6d3dDuCqyyebKtD0ClR612PA6jkkSj
pxyUMSX/4Rh6kJIFpzdJdOJhb3ohX3e6CG7eEVMGaTTVLgOlAuMU+gvtbKIIIwzVBWcIVfaQTy57
09cTldvR+ZUR03VS8ZHRjOJcarN2NLdGOwr0paAtUVSfcOB+q/AzloOvcHzNQqD3ybBykC61oO6o
HHFbJuUBFHkA8t5TkY7udnQ1IeUO1HZmATDUySWfJ8gm8LdzNOJVZKo3ivvlO9uBxBbyXytb9UfC
v8rwlMlecNkM+msHsmAaZ6vxPAgzr296rGBstJZfanHD+aduY9FWUNtitXBQ+Qt2ssEarjSUu3ib
uwmiWaRNlXKUtKXatRylIWlbz3hIz/jLo73hanGUfNlSb/gP5zK/EyRrGWTDnF6/ygpAEqsn94pj
AsibmW28wMJdoZYwuo1UyGNxoDerqjqgx/+lOUAs9HCXPxMAqCgn8uthIp8Rvc30kKGbWEFuh+P+
HOhrdGrA7A1WDHkESsTRrbx11hHng0GF7s6kIfHQi6Z6ywGvtGmYmIycSkQSBXAzArZOLtKSDE7T
4zMR1isS6hHAbRkbct2MqV9cZp3qP3+CF0kmTZ2l3BSSR54zKN+5Mmgnmk/FagjJB5kL+GiMJcX5
kc8iyJvIS/XeFurjO1exxsXc0/DQ0DhNUl8x6Z2eAv4r6tKntLoz4FeXGaWYfaoBuzhPYEzoflxX
ahoRYRyd+1sfwQosrvhn8yWXsSMC8w1ZVKtoN5etgxtFbIWfVzi5b/t+6VuvN9DyRrYyBNVpE8S6
JHPu6CDWsge9wRefJWhSVVxevk/1ha8OUwSmn6PPrwdx0t4HOxANuOyDdga7Z7/anQZkDi6+yOkU
m+X4fRPrOU1DdBdxQTZrrHxcfFlERKkZ0rStAxjjY/erYhNE53sxv+aq84OjC0DvXanuBY7kdPSb
VPHvZ+fnspHBOBp0VUT1h0UE39UxYUP9X0b1XU/jg4a5y3JejMGVyWdOFHj6ihbqlARhRu+hkaZk
epucKpRuoGXv/TpMB5UWvCGxqXgWkH8Jf/LhA9/1QSmlUsmbe/NK3y5EWsgc9YPOKeFJGPq+5cHz
jUv8sfmMhERU4l+KLC2C4/Wf/oPcj2QEq/lSaPKXNi2Z86gptVUQKSUYejz7RJlRdn+2xfqqQaN6
SSMArjV88YM+vcx42Z4ji4Pr8o8Xf74IVfpnA5n6k424piM/eUAUc2SazYJlPZ/isuUSYJ+bXlR2
OtdYgZQ4IHa72waYMrjwRo6hzdi0Y0cbzZl3sCCcmLEEGIbKAHc+VaPZ1SnTzBQOZRzIfjbJaTDZ
UoQEkPpNEu4OExVKQr+fS8ZvWgaPgkg3fQqxKPLjlZzSVjlydK5D6XszvN1L0VZfTcQDCtSNZPS/
by7UxkFeLrCkgO1CVTSYryzA5PFmhk0N+wHcvDEjw6Yt0dH2eBw48fYZYZeJVtuZq/8Hz91W5QJY
dIw1bnxJgVo+jflMxPQXHLPIYGHmi6EztIei7LNjSHtz3u55rceQKhRuqwvhuyAllVxtbszN0I8P
bKaHfnk8NkrCUdyju1NrizJE+BeZusOl+gYx0G4jLaCUeo08cFnGH6j1QgDcYSObQmlRPUyefxXW
XPQHTL2fgr1j6a/+BumeYOAXS7l+IJFq3nhNBlQRu/Xp/Cw1CU4OkGPavex0xnxBkEB+ldvxcbFb
LGcbd/3enwcubw6v3CWxEV60blXrpk2iwevCU6SSZBMpZfEX6EkVt2oBZ0RIAQkUs1dZHvs2IumJ
HEcwv5xNtygGuFb6fX5Xjxe8QGX4GnVUTvvgAOeLbc0lx5hljDugoF+/7w8PTDB9d6F0khg0TNs/
KmuVHmAWZk7H2yLnO76bWvC4jFzZ3PLi6kpgizRAFoudaAvjnd5Yqosvk/1BtYFsQnanzpWjmkqN
ADGRfTdzu82GbjmiRs9CKORf8hvah3eDZP1pq99Av78PDBtf2T+s1hqNna8brtLePAVcDpHJ9Ub4
ck3KNJ/5lunSk/HLnIExmW6fykn4PEAiuGjF34PtPCU8zi4D6MeuFQyP0o3CxQQzG8EDGMrtzbm7
nzgHYEeCgMlIGLUT41m1L/kv+VlvagBrFrsmOjHi4s3/vwTny5wE2aDrM2RRQPsXpJYsFIaEFkoZ
UFelFi8QXU4u/2GhkaX+Wsy7g4y6AS1GokLphVSP7YZJrTZKYqAUECZyYoXWKm0CItb0KvVRV7ML
RMNlNX4/yp4g59U1kbdU92y6YxQwH4w7EzZx92KoabmRvA/lVn7r4nv/boARtpEueWgqpjEdO3/M
Ezz1PtGbY4iFYG51CxdLkIdYyKDyASVJyr/EG8UJrXWFiNTo1HHPWLsJiO4YTGxOrcNZh+evvxp1
lXY9QftQH/0RqbXCniVL8M/mv9Suz3oxUmQ+RrouY6dykZomn0HbjAkLCtOl0l2LWiSotYYx2x+t
5s/b99BsBxJywATp/nOJI+ixpxPL7T1g0hhrBhqBaSE/At23sgPi1/IMJTXIzfA7ItGPErqhhT3G
u/PXq0C11IbAymqwfgWTPDWXN0LqyZhDmBs5x77aOy3vDaVAw0kRfAXL9voNfms88Xn74YWc6vAS
jtMBctT4+ri6edcqgSPhXzp7jGbfvN8rcbmrsbgywXTNyFUlKcGAjtkDdoIwpOyHKGpwCenT7Kc8
/Vgop2TxnpwvFePniDlM5UdvL6oRHqmUACexmqmJHIoiVa+HTXuPQbUbXS5i7COD25bOYKwc+xOq
KcrTI6HUPbSe4EPXZYrJXwQ+CfumFS75drkVLV9ge/my0pTWbS66wugYRYVtnvl3kyboFbFPafN1
MBPvvsX9hC49AIdQJz8EudEYWzfLzXgM/8OMyDPzFIQEGkJp1JI0c1ZQyT5G1GZcXzXeHD7JavBX
qVIZfZVZV4ZPFOsFKhI4wIkuqA0jGgrI4xIkN8zX/PNtELt4a/G9Iqn35qZuDu3abDjTyLvLWQAS
TP6u2o4pVZuSWftPdg324vA20a6UUPVx+Xc+h2Lln5acfr28w9rAVRjrEkcnKTcaZXuXikuYAhnT
oKdzpMkPHNAFwL/kvNrG2QdofM6Ld5GT/m8/dceErDJCTClEbJ9fSm/tMcw98hPue6xD0Cp1zfAw
Y0xlocqOqJaTYe1xM+1i0xomDTBTOH9ea2ZIUksTJqn7fDvFdg5m5GD+B6iIXqNK2DIkoX7EInjC
SjcIZm7dyIYrE2hOZ8ttB7WbgcOkRAHzDPz7w2FhSdPWDXrrqybmzoSz/7+EcMrMsnivVy/pYDHB
IlpyIoZz6rIXG4JHuTEox5K3o+8RqzlZawfcKFxquspwLKwNGmW5fX6FWMJ8jhnRuJMm5y5URWrU
zoA8xSRYgzYQfbR2psO4q/Vc114Vvd8V6liOuQpopyDcoSPu60W3rcn8A36LSM4cjrJYOkRPx/xF
LNtaZghRE9TARlyBfKazk2N/w0cvXHP6EeFKEHabGkEriPgPbWjaQ+wGxzS3pEh+WzGtt6ryeaPJ
HiIK4Nz4ZWppuAnsN9LfJRumhBJEmzzz8QpVZSOZFhQPz958yx/SLhhqyyIalO2+44sQbKT4vL9I
SlCb/c8uucWTp0KoogZ9KokZ4BRID66qMHvvDCjTTKY3+fAmKmPk3NiHIJRodEXtWQB4oT2M6lTE
v4T8w+WRZRKzI++7gkWVdBMjz6RxOfCTWNmWzS4o1dLR3rWMCgfYz2bpOpO37LcgFCsXblQESn7d
7Oit8M2HxmcN15HD94H5J2c1V5mFmWEwmQ+L1/MOh1RPpMUJuhpg84YILkp6x0FnG1EyGhHB7Goj
c/WZFcFs/SfHm7eebUjdXLylm6OC48QZDpyNI5tHEWLWLYRFdFcgWZIQoKL0BJRNcXNkDpRuyECN
Io/LZsfRttEFXksDPS5BJFEEpMGGtLhyP9I8UGCedhHcK5IKL/g4CI8Xw702NL0aEAAN4pCreV4Z
PBTgN9Bq4msE5vM19qzZ43uSI82MW1SIdau/wWsIysqZOjBPdp27Rnkt7KwJnxxh4yypyt1zMKtT
CcSMgN3kl6kxGbZ+0HadsEZzsJXu8V+k+uWg52WtJlt8kCUNSYh0A0DsdcCjufBauzMkMyJ20WVh
FpNU22ZYXVZ1MnwGtKGOyOYMyKHhH9aUWQuy0a0WOkhDmqsOYx2JoNMwulIT2Ex/kOaWTdpovj9h
cyXZf2TU13CxA5i8G76sKCtkQcJZZzCAk32m/oMPoehGXFedx4aTkhqqAH6lVO+zR3xAWPIRcXmD
DkeJ51W83YDcyIc+LJ8a3pKG6L9A032UFTD9TPT5m9DGHr1nwxH0b748UaFygOY65ahs/91YySXC
cIO3JE2Rr1s4MCyelOD2oGpPlxp4OH32yZ6PXRsAYCNDMd19nFX+eek7a/fKUDVL+dctEH1+oIN9
LFPe/xjGuqVvKcUhZgiEYSz8+mriQPYC46gWIgrnUhl3QPpjEQRd1lY5JA/W6jbWu05bAx3Kfnuv
z6t+a0zUaVBWv5NbwcTFCNQgerAUN3CLMJi9cmZrubghk+c2P1j2Gr/9D//SWfeJt1/NhrYrJ5je
ZOwcdgQHXVxaMmKM1GXNk0HOw2ciLDl62rPkQD+jvcERpD30fYZ5q5KOIHqMOxIJQdoLAi5h7wvm
AkywyE948TAw7SztaeOCMqBJNpXsyuKQr6DPbkxz4m37oCtDE27vVuWZ0z7hE4IHf+7q0gHEfRBS
Ir7ZxJbekqIsKEqHknbQXk//IZ1DbyXEcUI1cSxDz/r6feFmRyCl92BgOV92d7a8kuawTYJph6KI
Dy8hHH4h15EPHEtf9t6R8UeMFDxJtUirtEWMijapvzqkbyGqfY57eHA4rs+30pkk4t8BPNvGv/tq
KXIMKr0WGAIoX5wqFnT557NiSBRgUIW0RXmItRy95Ix66eTCsxcOyo5SScfTYN0ak5N9bN3game1
2OEvWC4L231M8pX1eZ4JK32as6/PyCHbH45N2YPnx00WrOFmbcOTKWrJ1ye7GapCndMftWOyLl5N
HHah3UiJEtAckglky0OtXa1A0KrDxi81TvCjM0ItOL0cMOZh6y24QvNL5vnfvwvii6OLWJNMp9Fy
DD3cbcZBMTVs6bDKy0TxirNXXxuGxuLcvckvSun7zVyhgQCH14KH+X+/KlF5RHslGpWJs9KgFpb0
DPIbMwHzwnf1jrK0hqwPsIn5SKtI4QWfiys3UoH5XFy5EOJYG5onv+LM7Ohao4n0enKxIaviyZBP
Mf+zrbUFZzxzpvJats96LTJ82/XxIFlrNZnwnZ4WxHRNwU94Pwg7r/3M+50IDavkGSFj+8tAkzZC
h1561i0nfpQEtCjatshssQ/DSB6r5rJ3bCAm6aDTjeXvvPMwrteKmN9KvJ3gPMjFBk0gGjw8Bihb
H547A4XvNsf1ADX1SsOZExcG57OZD85Zx8kmkIH3lZ/Ue1ynFmXKXEIQgrGITlOu6PGz2nUc2j0/
MTwq2zTVmubeXxZWfEM3ftUT1MxL2A1zH8h7MUgKNMSu/AR5BrjS+epTiCEN6QrJK5NPe9Tm/ilP
RDsVl4DmSv8Z4NlvoJg4QeyiBzQvVNyl9gu/nXYUxZlBJ1P1TyrZ0H8qXz44iAbqO3MXQxV52eXE
ZGisSa0PyxPnZ6N/v5WKtpt82CfPksFvPbz6y1YplB9MZlcv1JOBjIZTXL+hFqVsdAL9uFbV6uTb
NIJvmJcL+g3nx4nVv0L+KZ5LeWDI/fQJps2oorfReVdiFLPD1d9/3iPBooyi9VaPEv04giAX5S0F
YIS2+eKAJNvEGbgi39mi87ytjkkFVOtnk6Jc2QnGGvAhBywjXnvVWTXjSWupe4EjkwXxkNVgFZyn
iphCYUy+GdsBNe+/B2BZH1Pob3elbtSPZjgZclgi6dXW1KugA1Ah5OVKkogxWzOgGFPs7JFiBrMi
NLOAb9C/Z5yxa5U1Eh3GYnwR/WVYB8u8J64zALAvQDdMAS9vet/26pXZ6rsxi62RYXTWAg2lNzlf
gHDvQ/pOXjGa2HoMnHtJjB/avInLbSa62TmGtoejJ6J8G+j+B9YbN9BAvTRrp36f3DRRxLIkXmIh
SO/CIbgiloCL461GC7/k8DB3MOQlcHBxLtys5DZQL74Avi2k0JjIOBVv5VQalPiZxVo8aCDZ5a0O
HRtf4r/WTA44oDZxT6WJVDfZ4q4wcKVhlEkG7kSSEp5IHkJ+z1m3a99EUNEX/DldY2G/aKkp1Hdu
tvjQpAnvOW9CiIt4CTs+GtTRowZ6wGuw5Ge7BvP18sruCBYFjpKkZivmoInYDW139yvCntL86JTn
0MRDtKbsNOdQlzxvx5fVdV1RrQk+b3RGO+UTCZUnktvI0haf2/TgKfv+/ecdUQMnrhmqi2HY+Z/9
/z3hyElOX7wMTm+JJtyDEZhkwZlSvqwZWadCgKD88ip+ibqoeBNuVaWXfGMCqvCPCi6yK6ArIU+d
49NdUAk9jYxtxtuvFkKIUJpZOOHOl5nBefhCe5bnH46yF/lr3qt1tyk8TRw53Ro5kFeNZxSfWisT
qez5tvz9MutRYKYH8jYBPsrP7hL2Om/La1dMsCBI4O7Ua3ZmJcTSrzFL2g9MP8dCGdbcJD5Hai7y
4LDjI1ibbcO8Kxa4rw7j6PRZj03+bBACwpbtvUt/5v8gVrBOCLMVj3zFX+WYaW/hyyhRtw+PlbWZ
/MM7aZsiV4SJ/j13eEfnYbQm65DFLnxOjhLuTaf0AGiTDbnGvqwE4UgF9Y6cQo/IqaP9mEExdJBN
NT0pFzUpcuwIZ0Dc1Fk3C7bjl8vaWw4Z+DGRtoGjETm7LUMwRrJOSbewYCdFadcy9Jng8Pc44IOC
35lSYsVLMvUrvWKcIxAR2iL/hPuaCMv0yvWor1XI/67uyEBC/OU+ztJNXKkusb0NMA0deJ3Xb3uS
cVIGfWUM+QKYKofocOZFcj5ckzPNw5l0c60Xm5a+wNKAe69eBdknx9AxxCD4il6xxmuTDCOMPbDv
hcL4kAK6lJ9CJ4rcPLqQBynw8pbdHFYgZVJy7HSkgDy8PSmTsMVdmuMyFDjo5ou1kue7HboeyaRz
FBqFvvaSFP48LVN/cXAnJNqFAPz5umE6sAaSy+E3shojdXfSh1HEm8awwrj+Brur57tgnxM0csE2
+RQt2ugET+W3XdFXzNvRurKpIZM7VKbMAGWzhbuXo7N0FKp+7BBXSMjI9XrtwQTrMe1fNoX4mnHQ
ITf1gLAxNRVcULJZtp9uHZ/Gd7rugGgum9flT/GSq4zQ/kdWWNPc33ioGIUk4ZimSYF5hwGOsoFk
wwS136l/waOOE1Z5ltkkuHNkL4xWGouOE+szQspkaXdFXAv5mRl5YZXdpO9ahKYCv08+4oUYQmIv
tpbX11BbTeZPQkS1vOuE4v6x54R2QjtMqHASd2u7076hzowbFbqdW8uXshkE2STRBlb/7qpSUHbV
3udqSRv8xgmBq6B0d2AMNdZ5lSSzhhBcClswvQKi7vAXieoVLxKhgPJQ8lhacch5RryivLRkqcW1
R34f6KtCVWMR2anfTlYdMzuXaRlu3Or2+pVclvQsJVEJN5hKtkzVXfGc19pTOLSVAutdJGHMM3Ot
vM4Gy6nqN6lIm0qqihMNwRO7gvPRyX0vRrNHGZ6N5oMayMRngnX7tbCRWadeVmHPQiFSU1S0NWWk
r/c7h7mQgwXTutx7IwnZyGZi2ceFZLc2ywZjQHAoR31/dpfP2YEyaP0QYGFknS4tm8eKGd0yKFsN
7fk/ZGJIraKzPhH8iiC7cWYTSWzm7GNNyyl1ydU33mLXGYnW7Sb/1U2M/dqfR0zWeidq9wf99xon
UWVjWKZKyX3ITbzoOG9RzkZ4/BU6oCkFO6W+R0C/uaUFYWnJiRrx6z6EYMnqkzkyqiV2rSlno8yr
0QF54T8gx9M0MVDIjGuwhcEWbYjjcBW1DttDCCLLaitPcRhJw7uK12veWARERZcAnyBa7SJiDyMB
jTFUGWJcfCvjb3QF97Bc4dH8Ju2LMbaLgIYAcUTm53rsfKR5XPCqNPrZytpxOXYhlHG/tpobRwT/
IE6jX6km4kIuGvITSsKRtHeGPWHNLyZsKHrU+WBFCIZtXS5q8XCfI3zM5QRxYUPontJWwatxax+j
ZiU22THfx2HOPizooYLjdgB4PTOftPUe3T3GVNeEFgFMane8CptJY5/Cea/Mtgj2WXiG1WW9Pkgr
aICjzzavHc/3v4msZ2C4po7LqRm2mTwngTVIvijiTap8uoJO7kMDmazoQLsEaTnZ4BfjmlV+zymm
Scszhk7onj/CMGzVGSaMI9q4MASsjwYYm6YGP4AOmW5RXexawqHR/0f8wKJ+UlZ8edLCKsWPNJov
YMB/r4jqLwgsiASg87fz+JmfmYnYGEV466oWdufsEAgiuYcwpZiWm8wg/0EkSvTdn1d9yv+fhcRb
ZOPo2Ek6qMVd7PDNoDz02nV2l2TTuGnWNFU24RRrZGHqkNS+m46axuihF+/LIUHLCi4sLUCquXfC
5nDY2rsod4km87ECQsUiBHwMFfXcOMgofi5Cf4DY/HQ1h1DSojB+oJtOUSVCxXC0I3+AGa6xjpmr
H9I8MjNrXFVK8ohYDiYKgRqZSBZIc+tVZkd8oG/XaOlkOBkbpcrsYXJdxb0Mz8rgUgGH/3gU79Mg
pwyN68DOGk5i61Y9LTGBgaVdtRi7KeXbROq5hW1iVQ0iKW8G4fmJhs/o4nLJ4sHFbokiyYrm2eTZ
hXp8hYzKVVXCH6M7baxng1fwo39QYqMtNphCTf1GE8Y2FHtsTuJszpIbsnnsPqjc3l9QXMLemuXW
e1I+Y+lKI2kjsUsGejLH/FzRgxNWzD/S04sm0A2J7E3RRtsXbBdganIVe3hQmhowyGV50ooCFKZ6
qg1Hg8YiddOGIX21AojXjL6AY+xyimys46rDfIcz1U5MC52bmzs2XASqy/+MZzMkLRCadPLbMipX
vdhgac7WuEErqqPX1LyuObxE5sD9TZhnfJ/so6aMSnoXUfmmqiw1rm4+TMPxQKGmGt7NTjer0MQS
VphhVO9hHg1RHdrrSFPOVBWNZuRt8broBF94qe659YbtGg9ybY7rqD4vUhdDQsd3RtMPIK/nWEn0
t/zp1erh+MoKcczgRraFig9/z+MwyO+H1A8B3UbbdodtB3tKLNx2jRCHxViM9jEFLhSrnXRPaMdw
2HmwX7RfCiYt0ROhiLZkEVBHrWfgk4C4cdOUHbUQk5EOUq4kHXlMwRzP5e8VW5LABkDgK8KZF5pi
L8EXfwKrgESBpzMkK/YTL2HxtVHmzfUuULtagV9XeL48PNBJ6q4Jljzc+pCy+r1s7vYFVZgjj2NA
A0Moqlao3Kd6aqStbH6CsVMppHblp1oYjb1AILpdcLYSr2a9WFwBi/furWjYsK6AhAXYyWD2iMIb
RjCLJvLUUNphbvUPnB+1WiB5Mb/ppl3I3RXmqjQJEa5Jm/ESnNWEnFpc9Hc7cMkt1Ua2E9xrB9Qw
YA2FseoxU6PosHjey7pIkrpje3pa8cOCrrENQJmNyWr3qFTLM9jamfHUrBgNJ27HvQiqRCgO14ec
y8B2TrP53Hlu1UDLZLWADTAm+JsCAtJNWkYcWxV5CAobAlAXZROy08K2yn9pjt3o/RNAAGYhxAyy
p7hdSZq7mKtprJzXeoq/UWqvtJGzPgJGIxK8prMGILr8AgjHYJZBnphzghmE2VHcFeS0B2+jMEYQ
i2jKlcuZh7sCPOCS9ldmcQopbYrsEbeJDRYj4mlzJ4aUZIJ1hHpuV8ZYCqtrUJbNIeYev1D2RevS
91zO94OjXmliTVo8lzGiirhf1gxdg60c8Vk3BDmDRVWfa7rFAHYETlvHjtzFZpv9iJeioELxWjNK
6ZjleyrijdSgG1UxtToGaYuPwqQvGAHkyPk26eVhgbUFb8bPrsq825xPHbtjSxCQAQuSBRwLrMog
S0M6XuJiXcI+JNqRT3v2o3AujE8kyh9qzbMXZQxitQKnjVFJnzGGztf95Xj8I0DvyS6ONk+yb3aD
AiLjboKfzx7pkQqFs7oU8mWkmfpgCjGfhEr61IHg8fCocH+hmf93v68Qoz6rgK4NeA9xSzCyd81A
DYb2vfIXiBYxrEHkXUL2ftz6s7ZVJQgP4ed+ccT8ysxvD9/+hb/O4jiomrGGyHFMWPeGSHdKBpAe
SwO+j7p1ZDzvuV3zO9+aZEkrZhLbgPQ7L54VjI/Y9P1kqnL3SiIV1lkvhjJ46mnEt8Ztb6dGmOME
QtbFHoCjgB9v/7AaTyuFwE1+8qGSOb2n1fWDWZloReu7ElvsxLPQM0k8waBaGx6GwRZUHufjrik0
OKvLF0tSvRahPm+6qI0m9dMm4++IClh7vlbtt+ZVPjP13gAN+aXyotmBSF57h3zrHhfgh90R5i7J
tlYssZyk30qF2DKJv/Fti9rr8ZNnil/UjqiAPITc7hgbCvzI/9FvETreG2Cj8XPcZtulGRrrn6K1
7xZoZoIblE8gQ3NI0f6GBn3AvtYBh8uStyy6AJO9j0bnjX291hHBf0Bd+rJAWrYBn5lUIXb0Y6+w
23Dkkdw3lyIC0uUKJocHmV6GLI6u9byIrmNx52dRRMTNTV7aRtrl4WBV/JJIigSpjAiuKFSF5mA4
k76UcjXOHYPClrJ2dd2xb/4dI3LCDOvbnBYRHy41QXMKgrYf6B/3dVxsL0sEJ1/vQ4GHwR3M8FVr
wv/YmaOi3KSFFbODx75ymXGNA+EVgeUs7KPDWByGP86M9jzfWWK3X4PVCUrYGvD/fgAA8lJwyvGu
7uph8VyT/bOwflBBKc0SSlVoImFoj2H9pMvOoz6ScvJEX3PlY7HYtE1lX1JGPFfVFDBtd5+SSMnA
x59Hz3lnBsjNrQ7+YbClYxotNtVsfze0SyNBGiAp395AIH7I5u4wNuHxg6+vdpbEFtgqhIWNy2JB
6P47zcE7qlJEZ4UAxJBGt/4j1XtwCU1UGxetkmZRXlYJfF8Ek++lI9afMAt1iD6GcBXzMYkpGVHM
qYzqd1Nxv7AeCBvtQC2DA1kUqUtvKBlYTn/Cciy/lFQ5v70UvHjxmAPiK0Slv8VubN/ZKOfe88GI
G2OoJmau+CFeibzGuZD/RK/ph9C/+gys9um1v8mfIMLjYhVSH1JMgh5zcUIPyyrQ8ipTWbR6/L3K
bKz8mFqt+SDsAWvYi5V6wLxw2d8aEwYIkpMH+qqARuHkMC8MuJAaKqzPZQGJHhMstxeDMlZaBGZj
Hl6P/iUpyllFsIj2IZlZJVtwCXMjiiGHZIQq2/phDZRW8FqA741VSFYSMDlmidtqbxlYjvAD0Hbo
lYxcZnvJPAMg3lCk7bsBxSyxe34GXCJZ2+ArKV/91TB3F7+1IcXlns21QDacDTTDE+pnpXsyOBl8
RHTaG93oa7Bd745RtHTeRz6+uIVAkrhTQb09NubbcK6AF+9JafGNA0gkXe+LPIGIoCGKuKLuwCNK
AoJuZnbteMXUuyP9jxq0gmdnezBtng9pjIWt7q1y5Xrxj+vjwTzNL/WSkxpS8Ypd+T/D5zhbwH1m
Du2Uw0z5sJMYXZNSYuWW7mtwimvC/oJZkgJ1JAQOQJnBUoIyLBwR6A1/s0Cxq+HRiVDgdSfBDF+F
EjckF78KXIB5TCut61lnUd6ZNGFZ6Bj+SpUoU+Pn+sHRsXux7VFvOSyAFOjuFmw2Ik1R96opmw64
t5OkI4WvVTSeyr8Kmqhgrkd4tvnM+0QMezT8WAKd+GjbEKju028hZbSoMVzcErRPkFkOd45G9Tru
ynDOzZuwXZiVg/7aaxlgaZy4a1ze8xwaXxcZlxT4mkBfxC9EXSCg0mTfTvzLI/itHEgKNmlejFvm
JzRV0fbz5uxlWyUFT7eDcm5tbNvBocTgiZ9SHtuhoKAc6RaNuNtg9ENqZdcKa49jjsYlKDrJ3ANk
DAjuM6hH661cfUWpVOQw4WrdZND+seBfAH5bzAEGOfkPtNWBZ2UwCxTm6Y5AEd8MYwJcyxMEtRhN
ExGpbI/TroyYpauM8zcMgJd6A6y1X00n9RzrWnXJIjfXqbP8m88k8VCNlyacqRhHPoy15LTojCOX
Sn/zu8WDeejnKLkbf4YzOdAqktjXSIETL5NPZcYTP6jCjd3KflrTv4wVDWmi6qc8nCuw6mogglIu
vn8MRHABQwain2Jd1oyXAM2gLjxhPP4Oz3CJVZ8KV5m32GsobRoK5ys0rxEXGaEUnnJqtZNFonen
gEbdFtM5vFKVqATFkQOsrzRtc3sTNQdru/o2UMsJdQa/go+SLt9bkTeDp6hn4IwCZDHtKCYsQvo+
q9rMI3KEOQiie4ihHXtQto8W5hM2/m9o6IVjIY2bf14w1L+55DWWYN6D5Uo197x95NqqYPwgP1+7
hnN4T+yEaDF7D0SerCFCaD3g+46aSq7vdoSPafSscZVi/LZwOQd04gWTTLpHoYia5i0u5wB3YJnH
DNr9+rBB8G6v+1IeBMpNTFrRJgdlTbBiLlXeU8JG5rgOwDCs9sn+/3Rq5QD7UAyE4DK28LFG9ooY
e5SDbazjzR1OHMegoSpxh9WsnjSSem+PXii/jU6zYek2wwSdBgB5PYgPR0KXFSn2/mzDpRjuk3cs
x46M5RyyzcZyuc+uJz8oiOU03ZvD4jqGLyVHI+lym6Lsj8oc/E0PLRLt2pbMstItTxkZO7X5IDVw
UACrnKYVYD3gmk7cmkdvy51AmTB+lyB71uPnwHNuiH+n/Ef1ZJ2KIYqSwsg5rzeootXFaOwAsGWB
cZ7Yk3nEpsl1Bx2TmhAWF0xJ2zk6ET5cO/lJMcbQe8Fm85qMaGRYpw33j9iJWeIWTFXsIpNMJlJu
OD3oStMznAFtitTVuzNmDTZ6ra1bCDpR5biUy+sFN4rqY8wXnrr935VYeZQlkGHUdiKSX5knG5h1
CWUM+3sLGdtKICkf9IlW2g81FnvoQ70hhFk4BhgLMg1pqhoh9mzBx4LJZQf70sE4FY2YLZK+BZXj
6YB+HfkQlzBd70hu4u93Lau6Ry/LI5s5cx/74hAKw8CwhrBjq9/n4Ddeu2Ez5MDqAVGhBAciM4Dq
j7u1+MIgvfpTV8bdkeV7Mss8/k+1v0bJcPg7euFnRPX4ciFPXXcdIyeWtCK6PJuGyk1CJEJ69Wb4
CxUttBH+tlO2oGUcYf9wc5K5YvzSi+ni/fJtazu2bb27j2u6aNLb92oWggZTCKy7SdpeTL3cqK5p
9ib9wPLKNtv6eqSqIrGBSz4hIFKl5gX0zdPXO0aNtLH2VqVm8msxSizYf+tP4qIIP5R5mgmYsPXN
m+xEvs2m8g8kLN3czQNoB2JK443Li6mqFaPbA8FEKcrvWHvzCgXPLml0wVJ4Y5aecAr0JEcI06zB
a2zbiFyOAsHgU0kk7Wys/avO31ZGXl28HueaVJx1MLxAX2jI7E56uSghtWWE5j+eRzET16cF6tWg
tQxUdfB4JiZqwxEHEJdwwlepl8iOb4rpix8FVCIv6+BgqAQpE+8sM9yJ5AUexmsMGXLcly4FSLN7
bCB+JqIh5NO0q5WkRYS65kPaygxLdhnnuSNPcTex6Ebxt31ikQEDyxW7Mt0yTogIjgTXdrLFDYcC
vJ1yIE8uU8z0ixvxXdgJhWFQCF3YwUqw5cveZ8OzMLThyWjLEQ1AZEews5HYwDDHkemSiKxl4x5j
vhyaE1wyIJZsVzUH8WPD+MMDByGLcgoRXZR8b2NMnd5eg8hLP2G3Cfzjt0FFn25+wvPKFnd0mfte
yUQUJjXQ5XTwxv7SdQKNjbqJ2Roe527tirfU50mEyRAwExqFD71FIeDUvk31s4e+QiuvzNBeEMMB
J+kp5lVzfd67yKjVNwoWgHdPzagf6pajkPeRUvGV0ssDRhRBL78uej7UP0afCI+96DzRAK90XfLK
GSWaq58sZsRZYZRfv6IhL9XwqiMu0u6Zn1fdiM/3sZ5dZawJkSvASnJFD+Y1x7VUFRgPAsTLJqMQ
+HEGgexA+KzqyF8u2OH9+qZfK/gZmFHvLlNt/3MrEwBUKLgH/MTC1BU7jjR0juwDEGcSQItke2ZZ
Glwo4GwI/iqsTbMLWudCG3NyF7GWc+Loji3bEUNK5jEXbLyOOZ8OKAX89ErlPPKHXk1R+CRR56jI
9m+aCrJZ5Rn+581FFCqYaQjEHohpKe05HK1v3GIJDMNOztONlyP6OnbFwFq5MGUEe+UsD/NQZAVs
owSlhj8f92D6QGn6NmodjAEUB0myGMF/1C4AZ8Ylkguu4SR/NU3tW/rwlVCpHKJbIkIzMumNFZ8G
tEznC2iM1pSLSNR7tx+r5nI494JLrnEGwmeQ9fcLm2QurQ/j7pE/QCD3Vj925gKl2wJdkwW68VY3
uamoDXACrzztx1rnVqGMauHqSP7WQv0SU4h6Xv7Qp+2k3qsJSzzMeGx9jrowN9ZhHmc2I6ZsIEHi
LBBAV8vmpM3fmwkizyRhblFxoYni6UvdiDBS+eQLQ/83zz3YhOjx804mFUimansjbMb2zCnCu9GI
a7EQ2VQro51ve8r9mykEuc189Xw7L/rlAG5k+Qk5ypCUl+8AsNLI1C4Qo7w33DjEkc74GFW3BOzM
VgL34bkrO0qR+NxG+AOtMvmeiwIBw55YB+Y/AdWa3gI6szcBH6or85kowKAx8g2EFCOL99WU7zvp
kdmT63x4y75JwjqYJEg+PKrbbN6yvj4crTM8YR6rOFMys00ia5VFJrgn0fsHZLD5VIgBImDXiwuk
iRsRJapJLEbtntnZI1nzjBF98LuoU448C8tMrjz3Bq29qoEwkAQ7Kx1RD5Eeru/mlT5oaua87k0k
Wx+QHEyEX3Xjr6X6KB4/61RPmKH8ED6y/cWBUT4XQiYJkSXM4BauAd/4B4bWdUUrZZl8Y/loW9n6
KXIsfFMFTeQ5SK5WOKncK/wsyJqTqKOoOXxTff+IlhJHE2Km4UdFCgvSXTJ9rPitIPQO3znkJ1HK
g+SxLDmEMNMQad7uV4zNtZ2SEIN/Gnnk1T1G7rkxUJX6YIRpKgEYf5MGy/zVY3ZZV9w4VIr+ubvz
gkPqhhtZ3FlPaKIJoed1LXChsugNSy3pvbM5LFOpFfaF+wbdxW9JLJ/v9igcBfmRcHX+zeg7h8qx
2XGkQU+53ij4JLl/1TOuvVQ9GCopxW/7nyL1RgoLS5j16/nvbWQEc1W8vOlpDbR54q4DB4Fdyh8a
rOPd/Ays1Y9srtqrnGCL8Q0VjWuV+Y1mnlKg2O2LU1s+kDNZW4T34TJnYS/JBVaCVmSbQEGfIT/k
TrNhNJyttQVE8LuMEPDfjGFz3/jjWchpcKvznAbqT8pn4ET63mkkZMYz0gd+uHmYTcbxh4yJWz5W
zkilozqLYMv+75clTTU7vv1MgR7l6jc1DViynjtcWZJBEWWfoQ5VgntJnOXeeaibQhKpeXErG7SZ
iRb3/OKmqpxtnj7DXyY/AzTj+ncsN6NS1B+ulvCA20TEfaSWo31g+Dhc1bULY2cQLXvFxKMC/eOs
zLwjyfSu3VdfiuYSq//MlGMEj/+tRf6xQ9dkDMDm5fcdC+dp6Wb7YS1XIr4wuUl9yFgrhA/YPLVm
8KdXYK85HsxsFL90zTpB5oslQAmHmSZcg04SwvDMUFrZPpNWwXQaMdYszWszwCN7a4qfTZXIMpg1
1EsYxG7Ds8k0fZUPVzYJ+WsqwtFt3aSbivShSntraUeJYAx2SKzMwM4sSXhB+uzTHdxqfZx1+etI
7hL3gq753pqzm1W79+3n+qb59StFPEdf7DpG+KAls0Y3xv7hPf6jZiQlctfvGwq/IK8l+MQMqxH8
2cprUFD1ZJft2MVW9SP3o2FCnAQU5bzRqPklsiqSAOcGE/Oh8Rb3bzMexVeYrJ52bTZ9puI+re73
YTPbFcJ7XPLPeAZ2mI4iAtc27Wh8BHQAj9TowoSMKfPbnTjkRJi+W8idELjs4FE/zCkyQxEXVxWK
Ci1VYWx7kaivPy/vAtWpYVtfNbM+jR0sN0Jb3iQSsFsQIZ0AKYuSF/MMvULevofM+/mRXgpvIpsT
r5H1e2dxGC/qnr1PG1fUiddiZZcvxADKfsUoBDhNN9Wle+I7J8Dsb3iFYqbg9CaYH40/g4s6abfH
Pze9b2ze4V+xcglcsEalnPPI3ncv6mA5YbrrFrwt9KAbCLZ2+Z43aSJXWum6JBuzNDDuWdyQiqSp
x+pSpVWWwNVpNSQwlYft+tCbQ8PwjtO4R/jruaSf6n1761YrM9jLbm/F89EzB5xjgrZN9VaIKyTS
AtYYCVuCcpl82ZipG3iV/0sZtm1qgeCB5z65pc0mdSXyfnXWvcn931UJcVNzZPKAJVe/pdA9lYVq
hkiyhhh1qbtFBzIUhI9NtQNoUxTfdu02SOxya7luLPxv8H0VBvqNKFelCIiPfsX5ptLTuTc7IN42
nFibA46u+OSUrEGNuDP1O5DiUA1Zxoj99/gI1Hg5xdb3571fb4Sf7HGDdSGddwQoMUlam4BFL+c4
EeVEVmxnOrhl76601NTeIhbmascDE4ik718HrQW7u+nz+U9v8mtOErrmp+iHUdJSwU6zr6+EsmDj
JK0f1SHGKcfHB+lVKwXqKS9TRDZLj7BKcek32+LfvxxeI2BuBZF+gD4jaYcQX1Kh+obENzbtr5VB
8MdyljqOkQxDEUE1UiJMIvEMGSseufajVBqHkSY12TIXz3ep9QG357uhOJbPsX30cxX6sVKssRPG
20uE09Zsaq0F8/L6nmFKYTmaFBOhs6M7zAYw9FJTIaH0Dse3uvTPpuCE7MNnKhuV2oF6dkP4/709
PJ+MLhXaln14Uxb2wiNsy0Ea0Mtc+s97bvLbFMRnWEYJAWofue7NqSwoz0jfhomUPI2oHjUdwrKv
9Bt+70BkeU05P6cHkbRyVcq/k8/ADJtos+2ckrpSEjeE5vmCiN6oUbT6XxEqJciMomCQivqCIDVx
NXiHN6tbfX1UrkHB1ea6F/R46jFa7Z1OXimkrFrBGB/as1hd4Nr+HGnRwr/KERM0eISr6RdT0OlO
DSogVMEm4SXE3qJKUMe08zZFpiHenFWD4Ob/IeFWqgQFe2UtFVBlu5ZRQLDGZZzwrPTD/7VnK9+2
Y0p1giznWCONilCxY5wwaSINMQ5qe+DWVpyN6g2EpRLjE6NXlykrzFyaniaiCstSDY3lRlg6GZTy
EgPfAa3TDI/5IHKWYOMmtZqgvxn27/D5moj7MDYWXXCHOxgd5WKGYZcXBplwK63D0oyVyYPWYRsW
hbp2qfcxH5ZfGwQMU+iEyMommZjrwnepvqWTc1pPM++DzTdjuY1aAaFBBDJfFY+hpyTmNwgM2njo
foUqs5yNIdb2R/dx9lu2jZPAhmZrwfmJwYEGxbnyas2AAcWG5YhDHM0Pt7YSG4KK2o4r9GzLGDVn
1quDpkjA8kL9YxFf3DaQdjArE3fJYKYJ8WXqn7LP6iAWvL82m9BRGgSdYBkam8MtcwLC+NJFg0si
bdnwg4k5GqKsVKhSYGrJcb4/dx2LbTuf+Y4A4+JL6cEmsuB9CE4rs3NkgUpFyV/H9KLyAitbtTTj
Eb5reG8yE13IzXC5zwfgzb7RaDV1usx/PNvDwnAFRAMJX5oOw/qRJY9QKaLVxL/3ev+hOnv5u2RZ
Ck3HVSZ75RPMOgdQFqJH9CBKj0s2U+Pz8fzd+pFAJjU3kbuq5LoIUiU1zdRvag1eNI3ScZHGz3i1
mdE7IYoMz9S6/P5H+fP2864y9VhteZ0P8lF1mqWdK0qSRgTVLZC0MT4snqSxl8Rf7axjzbc5B0er
3Qrz1h7ASH0SZGjy0unYdopOTBiUlccCkbrvyMX++fas0UuMo9DDsidI5hx77E8438Axusaua3z9
styr8l/hjt3xd5xiuCvtPTtaNB7HepH9LY0ebaqPm65TW4fio3RUBuPjd9cKz5mEJRcmDJJrUTIW
z9aVxD2C74SvVV59ChKVjx7hv7VuJMglIGQKNE4p7r1Lqla19TpQfMg3UBUPid/cdw3xkd6bI4LI
QYwLwUth9pQRa720Z6motg++uaujwfdhQsQoESYcXCm9ScYfi5RJtqY8cT/cnJhbNeUcmmrEmW46
WchvzE923UHeamb8mFSLYbPK3drqiOW+nTNIT+uhvK8xJuSrXj5aLFZKz2AsTuzPdTVYstmIESW2
0yYnFDackrkhsvkESnCIQvd/NlzsQidGA3Tg2sEmwFDc0lZDzhEDpbceQcnP+qCwt/3BWD7bPeSl
1Bvfsgh45KezsTKDjied8lqkMgf5i9xDjRhg3CkQ0MSoT5SK2FCFCKkfFEV1XLIy3dLe9l4Ynitt
wPITNAbTqD7qVsZepTo3ZbOqqDfcSUKXWHwNpWirz3pM2U8vYeJZmKJbgEtxWAVz3iaKzLVR7WFz
qS2TPMXvWuxfED67Ej5ZSdeAcQXzzAn8E4GsSHGAAg1e+ov/crne3eN3r8UCoAxb/eF5jkBHWMyk
WqFoyjc8nnLxGg1IPSbG0cWXQRF9pwfeQ9KN1ugdIi576wnni/QSnAz79s6Aov3TjXTrHXxGGlYI
1HZV/Nmq0oxZ+Y9U/RSf3C3OzpKwWvp7WPz+1WiTbzjcgzX1kQaU4GllRBxV82Z/rQUNly6NBbPw
dXQd5jCoxFDwXftKCGOJP9cvTI3yLdhnF+X3jdU3IIagZqnCCdqdMnFRsilk8swRojUXam1K8oP8
yNM86dNUAcR6JoC5X+YH3nK1LDsq8ZQQzeoBx9X1ClowT84q+a7dsCZaCluxO4wKIqNpBvB9an7t
Lb7WF8qdvdSH1QyGbN+CAIdQi1+j0sLJugScW2HLLe+cGVVE0BZ3BJQ8SaFgg275YmdfJxermukL
Nit+YXyXfStjo+AGwTDW8OtWt653A16blUUue1YdngXYlHcy1Qoc20vei8qZU7r2rnzXe1g5jD3o
Sf9oiEJLcyF+bf1RK2zN9YwmLJZXh8ti4W0kyujcGr8c3CKmymaDrY3Z62845IIk3Tk1nq2+fizi
EPjlv/aR0w2IhcGr3/flOs/qHsoIg321svn1amLzGiU5PN+YdStJEDfmghBTmI8lVX8gYalbIK+u
GVEXBvDDrAhdM8W63ZCbjHBypI0qTaKZ/NUlgPPlV6oGIGZAcFjeQF4WzbMaA31DT9dpZNtcn0h3
8fxci8EvulwJUVVgmDatM5vwM2TNj4+jxVv74EnlTZpUHneMakiH4YP7dfybTpeDZWYgk2xizERE
m9fspipVGLv7sZhRxNAMe1znjFScrk17H3aK5y+ujR75dOfHq4pAiAexeCAA1hCiHzLXTX0gFhku
1AEipIdPzzvIOfZQp4Rr3mjDdZ8BiFBDmLF3MQnoF5Qvk7lCfz7A+AMiEklCKx3MpxREXqHfCli8
zMsmqpWg06PUGchTyy+eAr4u1mZaiUG1UxjK3sT672TaNeeZToHl7FgX0hnomOYS4uMFhp8BlYsi
jaNhA3ijNAaL/VkdExiquNTggaCophRLRJdl41HoZU11cXLg+NZimfuQlQnaC7Bt+QvK6YLNMkm0
wAJomXIEPy6tXiTZQHfp2IpuB/uUb/4QN4J0HFIL8orpaTndR7EuYSHfG5EbDTOV6CyfIGsZEzus
NA2dim3Kok5co9hklL9ib7bCY1+d5M2vhjz1ZKXBJ/FTAWZOxxJY+N/MIED1/4QjndUUADdOXOHN
4ERLl+Sz2H07zgjS6kXhBVJz6JwXCmC99U6zGXSd52dHDEFX0Kx5ca7Cb4pxh4dCIunch1/Eza9i
94XTG5hdcZp5X1NiBLBVYKl9zdMYLWKUPSzAbgmdaCnouQ7TgOEJhinX6xylb4bAAgfcIB2cWeL2
NGGGuNx9jeSwVMo6My6LVUFDnIkb1qzrqqjBj1IzA0w0CVQIUChzZ4K+YUa2PXsx1VtYu65m6eZW
uJbim93YLH/+ZOIYZhwhM+qqLsx8IsMrk/3OTT3qJaSl8WLSPn4qvXAfiTuWerLbLqc86tp0vwFh
TxDaBRk/ziRz2pBrh3p3rUKu+zvTIVjuK6vDg4eOraLipgNMWffSOzXbGb+dGv6gaeUP8oFGpff9
aPCQaT3sqrnOurXF7p1AW8p7w4JwfKz4a9rESdWydKFr6LwaTh+wo1L/3Vq+MiMTipi7zgKmqMjL
LIFgrEMkcC5rj0q4e1wzaogbg/YIKsxgWyvV6j/I6bOzPQMV3UWFG42V++sMCmA/iQ0RtZPoGmXa
W/twdHHmQ9THYlFmp7GWfmwMiQJCB48YZ8FsOOr91zYGfV+zxGTTDDCsvA0/Zyc0EAmarWITYtId
G4IPxGvF6UvkMCG1CHcdbvanPaFocxSvI3u6uONuscy2F/3hKLt3+gzXcmNv9FtShOSzifJL7+Bi
g8MGmpz3+wpfCGzDmQCH+n1+HqiZggPsuGtE1KrVA9UoLeEKDc3wsSazHYM50DM+oklcMkYIZoW3
FJR2D97e7ahOQ8oivITVanBxqo+i8aN117hLrU+fmnrWvXO98vnKMIjUyNmUZk+2NcpcYrOxVoKF
nhZXSWK6iHJCKlVl8opg5AJS65s+aHfZ6QYZNLHOCv53NapgzJDtTzKihg+CqxoWhhfrNRH18ok6
ff+5NZjw+AV3QuEp4jCWElHrJ+5BRDC3jXc8H+IayuHkTOc4mcp9DAtkGvJM+wiL3hidR2KCGu4q
E3iqBH4UOosBCBP8lCcl3LrGQRswU98aNJzyHO4jZqNjNu0Fw6BHr5YtMAVevwt410WGUkfvFFql
5Y53MCngL1TCPkMHae2uJQJslyL4n7SVROoo01FyBKh1YINuV/5U8LLDVAiNYzRXSLvIwx4b9n5G
j3DDs54fKK3ZJ2JFeXM8iEZyoM1CAaiLYZrWcpwQK83eulUME08fIrm7PY0CEqA4DeuImsnn6Fpe
VpevcoAGanmauszpd3YAhM2ulbORvptn3nV1AFbGf4/C3NL46IKUgcUz5kTLUR5qXA4I0EsF/fOy
PN68rgUO0UraKdnfEQwhVMUVfdjulrV25CbxPD0x0PQIbxx1zfMSxNPota1w2XfksgpKi1wGTCbV
WkVhct2hRRL1lkiF0NWjNzn5c7KDT2rWiI1M4pcyPrcvPSEG+wdtJBzBaIVDRjuDDxKASPHpToJE
uD2h7lk8IamZ9kig9Wf2wXNu9UWr+6v+OGjQGdqPtqjS8XJpYKZa8qCDQDtWwATT8AE9U+q4Bj4K
gC8x2uxDB2X3v0L3BH+dZoQk8KCyn1lU/T1jH3oxMEukFpRTWImxA9/jsIdQVxpFup+Swo2tkfgV
yZGJmqzQPELwPlhWKPWB3Hs+fJQxnuJJQPlDi3S8c43AX0J3o0hMS2jIacVVBFMt+v6QMcXO83/G
rDiVIUWChpW51dUr7HMzHISwh6W5tYopqXrCEKRWhBwYFxyvxS9yqkKh1sAMDz4/GkacteSdgz4J
yh33hxRCmllz5+9qHfwLYO95uPpGiA6a28lmI9chZxChnlYqWIZEgMsEtOktFAKagSX43BeCJLa0
Prguhdv7HO6MeJlEWS9ljJCc2O+JE4thDKD+MLyRQ/H4KFFqvMY9f7EYInIql94pXhpaSFby1Hsm
VwWqCaCp9pCvfhTh+lNHOKOXaQfTp733rZoQIr7m+Ee/JD0aCzI1fMjZp2Eaa9Huh0FL7rt+UotL
wPMbhDrr6TwYDnRTbbKBlP74qUUsw1MUw2cm43ElSgeOCg3VtKzTZBu/18Wj+OBUF86/CL/jDuYk
AKiZLg/PllV+jprEwO4N1NPtYB+9CvODsPJAq1TmxjDoI7lugduWHYAENQ92/72OwWUwxLv1C8EK
XbgkcKkGYMujGKoG8JrFNWw7fTQeo3JwHzuDSrX9++mPTpSkp5HYpQJakz5cNjC1e0U32UoZjHkf
/r5PVPzx+ynF6DcmQylDC/zcRzMZq6PkeRM5lDEKYlOoHRNxZMFTiekEiT0LdDncGgNNaShoQsTj
Tm/oRksEcm/+K8HpXw2sJPBasy4E58ss2TBRYOjxmMOvKpmYAaO/dCpbVkz1deIaTJ3NJfizaIKW
LdXtUVNlSwo51GcJxWFsrTFD1l6OaKUHNCby4LzjDnhDEgrM67S1FMkOzUE5o4wk9sEcBEB03Ocg
1RapWVZbF9X0vQU3s2aL23OQXKeQK7o7Jy24iMf11fi0odGtKvxphfhkNhvAmhJFvdmyID3uA2R1
Iv/uzhPnP4wQIgyvvr9UPyW/hrKf9m/eiOjTV9EdgRbqr+YXv1xcQETaViw8DU0JuEbIjatJ1sCV
NKpOsU2jPE6Xr/CVtQmnS9IM2lCib2uN76hymVw5PLd5cYwx4c/ihvo1Msb0SOQcLom4/cHf/ztx
DW1eW7FwUpbGVJs2m69FftsiAmTAN6yqbXhzN/Uuoit9cZGpJxPJuKAy83V+C4S4WW9WN55M+uvw
Vr1XKZm2L7tKAtoKYqtQKek5xdsVnlU/qWicMa1XBBN4UqYrrerr1lZz5Nf92Xei0faY1Tk4JBz3
dqS1aV2TjKGl9CLBIGq3OC9n0rX8Rh5ynVv02Ci7JlO/qYef9NWPNlrQvz+OFx4HgZCB+PZY7laP
0xTjXEWhrbxKxMNFkGoXXhXQV3zYM0oBRLU1jV8JodGuw3WUjE5x90N7Ovcfjb9jU6Qs7K7VbFFq
i79qpJGB9WzUkcNh9Cl+wPAPnxR9X6wv0vUOm7HhC8tx5onNEgqSesVBQng4fIcdfxuM7D1IM1B1
pSRiRoZ35GkqCIuD9zH+Vq0I9ALI5+1SCKNVlYD+sPPQxs54wODEYbsLcl3MebteZ8ZA/d3YpEL6
YFlaNjsou4ETAWWMz/uC2tXoaI5Y0JmM29tedDQA3VM0eZ1AgqNDd4TWxeXxpOgo3x0x35gHxuZW
CIRIvpJ34RaaRMgLwlp+SBH3W+9GkPO1M5J9KIPvik/ovBpWQqNUCmEQWwUZ9/kmc7PQ184xasKd
AkHKzUPQJ1Tmh1OtPdjt5TJ2YNPLMdDSpO1mf/I+Czb47SH75QWwmY/2vVm8v93WH6vlfO+MRRUr
OLSRQUUiPL5Hy1NCQVi1gqw+6yfgdGrq+kAtVwvjL78RyRCMO3NT1xo3iTyjvRbTRWGfN5pFay1n
gn47IqTx7pMVnZedvVItbL7dLnwhx23AagEj+cc6aeBBDGAHSrjbROrtGHDE3rHuiAgFmT8eA2ip
Vgla1GccDFDFuQSnCECsJ6T99pZA3r0cSlTlED1uyedKdjzAev59duXEbE7AT137VR8uSW29xhAo
TIXgddavQvu2+Xmz4DRHirvOuIjNRuQJx4kBSHKc12wcDZDamCabVW+eaKVQDsOHwJQQTFOiYqE+
6cv1Orzbsxqi12W7hS883X8AFCMwKARVQXbn6tPGH8Qk77PJWnHoU8et676g1c/TQUx5RgDN8O8x
KE8YwBt7P+4GP2VceJU0sgXotS8ZZG0d5xgntiTC2qApMXbo3TQIlWQDLbc+ZH92zxsoTya85FbZ
MOY9PXjb6Iy6xATAB0tnvpF+sQpDFipANQj0s9erYe3tNqzYYZbp4ldGcOjOq2mCUUkDhyhhVQgs
3/4Sw5uWPiAuXNdD1M3fWOPPddc3fOaNism/xlFMR1X9Erw6bENEohgCHq0Ct9u9qCSXwfalzvtc
MVmtNP138U5oNUGGLYmMoZlrDVuG8OERs7TXuEdxWZS/vKwzogBidQOKJKvyWlPW4t8SJ1p+rx1r
YVwAFStzeXjmKBB1q7Lhf6wTLXIaq6bp2fx5zZCyYrbnMPKBsFxxWwP8t0Equ1BQlVN9lmX1DqUy
jmPwhI8Y4LEEAzhRSdB8OmYKfpEivg6Gc/PQkK8bipis5srAO33mTx10VH94OFN179y8gYcbB83t
mNaz7wpmGVy9gQZwooV/bmL4oQewi/dUXSFXYX/KK8Zj292hcsZJTMMopZ+M13fEej6X13I5JNHo
Oc5N1iUFQ0dWGdEeharfKnL7cDTcESk0ZkdvGKWFgwoyVrSYCKkodNOcUiweJprXpzau0LMr51OH
9EHBNgLSWFxgB8OG9VJozJG//F1ufRA8rTsQ9KuPazZVO9HazDONQnbq96iSUzW8RecKljKZeSIK
QumBbTdG41qQlhlnyObQXv3X5tlz5/f97ig4hPAE4LDZPoOODehgOH+J61nAlGnY5bKlXN5Ka/xs
U9yAgw2PwzECEA/msg6dn6jU7pyrPclZi7f1Uklnu/SQ/ZViP3UYgtqblmaM5FhCW/3rqQOkLBpf
U11+kYLaOmJA79H/4OJNuRlqs6yTpWL6MkSEW0GFl7v2AkZg51Ngg6rz8TO6RoU1lAk+jZ8xZNUE
VENRFhuXZK+95T3zCqfYa6XvVGvXcwheOScnyQZFx/UVV21X8vEBVRknqF8334LxiOM7ByuZV2FT
+uzN0l0aC6qzWTLtBUpVFaxsVZ6ORnuA7JXXODqxzHS/D1p9MXKt901AUdA11P8psWBokK5x1gQM
gd2gLyCOVnciGlJlWSelRj0cg2xLuGf2Ygg7tvUA8n38BkUwZNb/zl6WhhdIaS6SalZ9nwyds/5T
0oGWHrfqDn9aS6DRwfd9EUGsgOagGHVzkGiC0Czc07NgY/HNsDQ2wLty4iasN2Ht9hVaZi7dHthP
mQsDSlwSAcIOJbfEr0EAgGcJmu3Vxc7nBXVPieE6gM+yIfznCs04cbKZHrQVEkp0mpapLr+6vWgf
zeqwVpYTq2t4zemCxv4pgu171kfkWUmIXPPv6U+/zzmr/RlV+DSS7160SYMxRWcvceKIyIqz+MPD
E4IjS8nQnPW4XMd1pqtjKYqFHY5TW7poco1sYs5IlGpCFxsVuE1QI4H4ixbqH9+VLrw7rvEjt2fd
XsFg7sNIWt+cddWi1/bscgm+pN65ZiQkiLPrfwsqLOQRJuse5ObDohxDHcMglz/MoRG3O0qYtwhY
drrHfFL7e8QKlLlsJaYlcYK2s7d3PjDRzltQ8sSiddw6zlOPNrJnfSaMrfmdT1w9K2BS/+8khhnV
foDS7xgc3G1NEyG/xL+ct1kR/Cj2F6KtLgytSR95TjRLYJLhKiNSirowljJPie/0niGrp8Y+fwBo
ICaCsTPgsLOp7iPW2k+IZIVdkkMbOEyTl6EEatEROcC0jBiJxsxXVMUwMqU7rXyspJMOqzn2H100
tEZZZqSZyaOJJLACD4MbQqzHVpKlUiiyFtSRxabKg+Fb7+/dUNB8bguJscD/7f/a8l2YplhoX9xq
657LH3PjsnjIOgju1hYmTQJf4Y9dD4A4fI7hL0sYgScnCtjMqbtFwIZnSr1UvmzDhMyqr1CPFtme
UJf+G6WWhCGtEejJBsRkDZjmAyb4HSyOs+GV0HH0LAab9T7tG6f2/PjYnqUYwOeX/rnLxYGctDIt
LHoH1lzq/k1Yy8TUxocoXAebSYIu6FSe1coUvy1Y7lFLH4VB1FFin81rP0+X58Lniwsc9TEugBFg
6b6MXId+FKSsIOYgMdDiYBPrXwqCNyu9X7kJMW4ZPWMDaifqhKTnAJYw7aBKT0lM6TjWkwB+1nCC
NMe/7fHciAmo75vMw5y52IAsugOgDO4Ap2uhe0Wp3NB1CHY2trsRe0TMynZF6FeQe1hYlb6Z2bYX
N5HSkdjgbEltm2744gfalg2cU1k9OyK+vBw+Ns7jWUQsxer4xH9lb9AlWSYUyedtjI/JIv1sN018
LI8fPqojUGJErM+zaJ+0TCDKnHAjLQH7oyvXeCwGlTjRvPd8gEsKMmTonI14WFtiWWk9fyCxjOOK
cNtkrqmM+L7+DDppzeZ4w3jVM7ksP7j7cKEOIaMi/p1VhuexTrK40ipmcRDSw6B1jBdXNdAQcAwU
U0bCS0r5zQ2x/u8ulfS+2jIi7j0e39oddEftISv6uCnoetoB73SzCIdwQRnreR4bT18mizL99KpH
P2p3Yd2dL1betD1KQXHjPs/GaTyJi4gKLH9ao0q7+JOj6S27kQQCPp571SUrNIYBpdqnx7o1NBYm
YHIcONGMlzFbHWxHDqRLF4I1lJYanXqbJm81DRHxQIajZ/N3HPhQM7cmnAzmge2IMi6ACrjxzQdr
D6wVcnyejSWWWXEVmqO1IJxrS81l5f0mFzldO/W6S4O+cMxZn6Fb9o2gsLQrH8QdwR5VwVoAw5Tq
MUp+nGuRDIrEYhWqQfy19vXQyDq2UeAUuCfefJdeXkjc4sWlF8cuDWLpuYNbOBPcd3/xKcWAeUf2
xZatHqgGwmY/nWM8n7T1Y9CMWBtQuiXSq3lXlu5vq59/cKyisIv/F24whqpVIZNLEcSGHfir92+X
uXPW75gECigy4dOVOVYMgLDKqZNraZ9V0ve1eNDaEhFapcrOjVbX3C8NZRZnY9BLVSIsAlst3rQp
d6VWUCGLEIAeLYb81BOrcDkGGTqF4FUQ2YT8URvbQpfi/C94Cxc6vbA40JFaYjE1M6pLHpdmuOMV
Ob/YlcLpYRKaJ1I/ZGykBBCn0NFYy/6HHl6YRX1TuP3KapzgD6kKQEpDyxAJdXL47ultFogyuhw2
onWngfxMnd24/uC3hLvythUZwqjQUNCAgGsArLYlpZwccDYHyho6UsDJy5ZK7MyRAIMc2cQE7vP5
/5wSa0vcvg2nfT7qwIq1CqePcbUUOIr1LijF361rGoTV0R3yk9GvIMSFfZSkOZJ58zQ/dkOCArzO
tVDZQO9w/3EX2u0BwbwwtIqDALhP09odItGjjrKH65shA9xvEsS7rGOqPiJxWRETBBfOrZZMh5l8
7spIop2NNc0hL+DSVB9Hqk/bAXzrhLGBMRNMnTzWrHCCTCJOs59hMOVp6aTqtdgOCL1OM7G3pTeR
2UUHKUcDwtgcf13Ggl6vrLjv3MyGamvM35nE+W9Bg0cWZ8km1av2Ec9HCXgFgNBlcuH3wA10+OF5
hKBo6TcVebF92BslHE482XMGOWhusD8fs6Vt+xTRRpgCYHnOQqsLQ4bkD9g6yLXrpxoV/9qxSi2Q
tOcyD5fFyviornh1cmJ/piT95gWi6Z31ZlSyoWpyVWs2+Y7kVpcWyB24uPhUVRWgKE6eja0KXQu/
betXCX4PBsJGPg0C82du/mMsFcAj5GqAaXDM9bPhhq+PtuyVgwyqkVTCuHM8XZOebI/n6DGcneCh
HM4QwAsY+jo5NlrKnvUu97MZQh7GPD+9dW6r+/uURx8UriEK1NZPlpE/kk/FdKeZ9udftIgg51WR
l5PaTIRliy/Up32Qh1wrOUITrR70/ikGF3Zjkg2DK9c03M7LPnlrgEaB8b67V5U2QKsYK12OSj5j
hkZDoydHLB6lwAqFuczQ6E4ZGR1YPYLDTKbO+8EKw0b29qvkiLKDxT+NoDts179nIp0z3FsdIbs1
F30BVd3W91ICH3zU/tPoK9XeO4jGbY/4QRjTN0rhwYGooghMpXo+EMndG8UX32yIifrewfDMO/PX
Qy80IVe+AHYPq+VjPKMpgwSlFG9AIbgGrQtuOvxzAYTnFhjBsCz46rkAgwMtl9P3o1as0QF6e2Os
7JSGNiXY8vit7ggAVAifQlKUNKQSi27ku8Rx58vOSVNpCRjzTl0QfNRCCjlGeW3NQjCkyW3JvN+y
1Y5F11z6bkT22Jdz2Ptw6rE20ogNnoxMAyWH3NGsc0kELycC2BDFgn6XTz80cdFWKQbMeSmsAzGY
9q8iyU5m+0V7Zo+/CmFn5lrs/LkF0zAflYzALGItq4iGeDxOCv4N2eh9S26GAqWc3hcDzQluv4ty
UhdXgOMFrmmb19eaQyAXPQcKdbgYUnwJV0Qw1koQsA6rI5Rdh91TDus+4bhg77dYIeMSGMHCaOQG
muBRFq+FdIqT2yboozEpOhNphFnHTgv4LD1I98x1whD+YMKej0BNGGAqWeE1WTzXdBUl76+4qerZ
kDepOrZQWdzv+aDcVHMlGWvEk44jMxLrJIz0NjbNKAOdhrRnqIKcC5J9P+yk7+aiipCZlQ3yisdJ
xKOgRl4oYCuEjzfgh3tDPujehBcgjEr/zTBZYkxN9RHqorGLkn2oNhwcio5JUUQ1XRMjlR3fijzI
STX9s/lfcLN3Ngd9O1LDgFnCAYS18k44vcMiCWJpgJeXKHsJRkmhTMrOFy8CKw4fZiaKga2rRcFR
5Iq2Wekgmp7ZzzRCIKmvIt2EhxNNgg7BSGKh+OG/w0bLJZ3KJNCX+S2z73Wqrxz3puMe3TVCsVag
iO4osby9R/3XyyCMR8d5DjAi595UBiVkTUPqCVKcCynWqJR9fPWDBp6pN5izH5MhcACkrfZmEpvf
Y5yfjyroH6GBBbSmI7tk36oSkGvdMRMTD6gtqZaXXdftKDbtxsG0cO+1CSibNftz7qHuSHKO8mf+
oj7MOHm7PgAyh9ZNaceitwVDeNOcwneINZsJXQDpKlxjz1zO71djOPtctQzBQwU11ggWZICZNPZS
tuvqiMPc+u7FJTy9QZmlf0IxHH2yOqcrHPDVmALfZOIBMlkst0iDe2vn+Xkqo8v1MV1l1Y9M3CBm
+9HP7amh7db27sJPdXUWfrjDCJOeFfYtPn/6QB3z76XvnBvwGBHgua4rHjJoExuZIcBZ4+v6X9WK
jKgU+49MXMwJGWAoVT/UV48UE6sacM0rC7R8NXF2D6IXfJiRLYGKRHW/JIZM+ray8EkbYt3K0Rxb
zP2oEYKAQc63FiPFmOO49k/PLGPHwd1YX6ukmPUV8NM3iMhrcVdFl/RWKL9S6y31DgC35HXyxIF3
QJiCKknEZ80NRJgbBx+W54V9pGlwBuTzh6zoGZt7mKDYO0nRXhJSmSJNhsPWzPHPT+zyK2JlCECh
JizyZ5HF/YzrUpMiRPlxPwHJXUU9QkNfrIGFF9+FIDl//ln9Xs63DijHYdMCQNem/i1EJJ32qT08
qq3An8SVNCzkHoizPPEw2oJnVVVVydFQbFoZdf+sq6fc75aPQfpdF1H4ShxKuhaANZezmuPTz5U6
by0pzj0rnTZmcxkelbCGPZs5TLfMyKaYBMpsSmaTfGLdbJ6I/i+j31+qBzAzO6D/AKQ7fgvQCA1Y
8Oh2uDx4x9rAU96gZxqrbnagzaq6gNenvRvDoUgjaDAGEm7nL+/yF4qsWyAQHdsLuz4fbAuOmDaA
Yvy2MziiijqLMUcFkPRkw/Pwov7nrtk1QUFkESn7xQBjsPZjdTn8YXxRE2sbONXcGMkBK3NY3yfy
HV8E9tIfSqawUeE/a4Nk9yYxkTOhB721PTlOes46nSkoY/h3Ke9OAaVFZO4SWIpvL3lVXgV2eLO6
oj0DNlzGMaB88+V7THFxvsDuE2X39pyrtfn7ujuD+i1GOd23jrkO2Wn5Gz74+8fMWHoJ77/gcdSi
fANxsWtwZL6ItLrs+YfXTox49oyyuy+C8rtCKcR2nBH4M+7AjF9aODr9pzuPUo3jqISF6GzzPp/b
E9HjqBLJZhqEYwxczBUPk6YD190geKCi+HgbhCzyyZNwBWwI/ebQGNTgfYJ1eC0qCDY+OzkpBCKO
FY4+V9QL0pOaYy/UIXj6LOUtVtABVLt/oucRuQGK1R4/NKpc7W6wCcJsD9zp+PVvgiMzwGRubiRJ
kBP7VCIxKoMclaWAgGu9Jnc86G8FdwwawZCxb+BSyLMo/fyrMM4tpL6T5KbYbIGm6WuOe3pWykjO
gky4mg5wVr/u4EJuTnuX/CwhKh7+bTXaIGS6uS2zH0s5DoWw8T7ne4ytmGSsTUI80hq7fNTt/M18
2vQAuenfGJPQvYlSh6c8RhBXA7yaCgpr1q9KzA7K+AuBzLbyC78a/QNKwhXMlhGmoptwEHA2QtOe
NEz8Of6s/5k5RhPBO3Nj6oNl+AKA0fOlQqpzjFPCyIlxMvjEt1f30oUTCzGphbJ4e2FIlzhqrH2M
03Y5Pn9RuKj4jlVaR+blaFRtK8J2uAOo2bBDSG2PYHVkcHu4Cx829TSqvkD9Ib4bR3uz+HEIYnXb
I3+bEsvuPssHjP7B+wyHjmgmOcevQkTfnzRrwpLizTILf93smRX75Rah4z3wwtyxP7KXXtnG/ehn
2OTUt2eXpQx78d1cWvL28P0NcA3TxkRMUzNqtch4aM2vu4XG8BCy4s8r8ycl72HaktwWT2A0Fn4k
UlmVfiS2RwUrMfJvwMo5pP6IZqvyi3l/auu/K6ewqKys/CIjhbZHVeaaaj/azybLkXPpgTHb5TFY
0qIAxamnaAGNcOmj/XJY6f+i9RgwpS78OK4w6/p2VtIKSb2J38RHMyanmFTjGZ5VHwBFLZnDAfnj
BJq7TpLTvt5VSJM7IaYjJzsZlLuS3Vx+POaqIwWwiu672E+aQfKPUjMJKEiHbHAf+n7H3YHQTZpZ
f/ZIHHvRf8kh2JmyKpmrrf9mLZyNxHFtLOion+RoLA5w7U5qQXFpNoVnMTIZ8GzncmbpT5TE2U6E
/mxXon+xaMxsKhXsU4keBH9g/NC1cohLTMLcGDO558XOE++13tpgaIoG8JV5dOQZU6YHQWThNDUK
zmUkU2NZFH7RvinPMTJlMaAo+4yQRs891PN+pm2EJ3hzppBho0+ohssP0EtKQtK1B4qrh8HVtJn/
5ytrhGKwPH2BJwGoiFq6pD9eBZLdOVz7pLT1qbKRdrDhUILDaYFaEP3STNK1jBxxWApHYbFnx+eu
iD2ueLElBBGiCH0F6bYye46+sspH0ZFxfjocQ8DneLxs2TYaU7wyjVI07K25IYQJ95MO1hZcrDZK
MBBQn6K7YsBT1X4IRedbclzevrv6+FmpwgbVBk1sKEdU5rIOSKNMqlfAqpRLa8ugeGc8E875DSZg
3QBBI2OtiKywNRSQVp3a2iLTHi/SQPJA7B5DdX1eEiPq5C5ODmqTlzdYOytS42M+N+HXNAkdHMkR
thNCkyBh3O5LYKGpuVx/P0MPQKLzAEg93nOjgOP+aPpt55ZxZ8e6mi0ws0wjqOIB6RRtuMV0e8Jb
g0Xpf5nVpnhPFwSNEg5138gzjbxToizAt9f9R9qDe/KbLJAAFXOPAaRYdiJePF5/44GZ64a1e/7r
wNR1YV0qmdAuwpn1pJKfY9ZVvXttk61akHaeUA2Xk4iq1fNNK/oZq/OBefEoFCfkBmclZ7GuevnA
XnOHYMLF2YJDiVYJJLMya7FL9j7zTcknkdLeZ34o3zAXGwI7MvXQFdw9GHV3FLxicA4twQu3iRSp
T3KuhzgZTnrJMgifGZmtg8X+OgOEJUKSceLEVnfru0weU9z+qZ21Z/XT/rRAqvP+XBRwVD0vgTfA
CZxIKh4tnSkhmFXuTZdu1B5dLJ1ZWB6W/N00NqKBWlpu5AT0+Z4W1qbTMYiui6UHTChpRszuqqEw
8ziI2rModaIkSYTpA0hGeXU+O0tSx04asV9x55jSrxgl0tR9jntRQSkgcsNI2hIZXDNEeo4x+Zgj
gMRvkmNwhXvGHLOwlutBQoBYrZqdpaqKVNZVfYABQh1smoGJ/mw0/dCgBih/JONgIX08JV/SzW6u
v0l39RkEFmh0mFbaZ4ZiUe/oGx5lMqiWR6hkHM5tcjf7EhhAxLZd191dhdoFxsL3TvS6cgPlAfSL
17ec5IpEJAesrwEW82uYrRw2GMuwEvf4GVo6c67d0QPD5WPhgxPsaIF3HL+DGg9L7p9t8sw1VcNf
IWXWR+Y6wV3oLEr2S/CHsk6MrfJuZZFDxrfJ2lj5Fc/G+WkqpJWxsm4jScFJeuj1Ys/wXLU4KdLz
Tu578KzHVXM28Mu2/uL+p6l4TJwDm6KgVaE24orzyF5rcgBfwgDFcg7cPpCeKUwYXSBPz/TtrIWx
Lvtd1n6x03boTA5BUd35pyCPDOiNdO/vZMcyzNsU9dMy3+TmR+IWS3JTZR3v+pvocV8r4on7q1SM
z6rjWotIBd9RKLLGeZx+9gtpKOBCKEPOZPFwTbbjxp9JBMMBDmYjvEF1u4sRHSH0WOq3Td6fF+K9
u5bdG4NMthMC2+eqy/YL99OmTxRA8KERDv89pje3i0GhgGXuCZZPzoiAPa/qOnIWhv8+0y/vbh/u
B4Miu6RtNsuulMLbeB3b4ljtVAYcmHqubg91hOcSkXivUk8fCW/W0divLvzC+4eBXWZ8xVu7ebrV
8ec3cNQ0ekhEMAwBR47Ef8BUYlPAgXtcupDo39qvWojtPi7OiRKt2SLE0x9YWRRaERo20uPuSdIg
GRMrvbOHauv+qlelADy2ZD2UlTr3N931CrI3Fm7XDadCSMYSZdRafnUAIeKloU6jJsl1lQItQoSB
9WCDALTz8IWcR+hQ6ZXdsdgOTYTMi2gV2vAQtgCz1wzlcexzrvWkAcjYs1Wxh8fjJkNROg9rU5Y6
pttBWqqF+c63ijglJlHwNCBwb9KtckS9x1UJsZa59N4ury4BpNFbCjZxCXOxYv++VAG6rLAn3p7X
IM0QVPeOyqYpj5KSzaj9Zts2vido/khSZCXHPliPrSQvYfL3AUK2p2XsfxS8sgtdM9Xbap5JhU8z
ABKCE3Y0lUVPwrwiPDX/8MgS4rHa/A9geHEd9BtXLzRTdzT8hKmFXCZN/ORPW1QcXIBC1euaVZ5I
KakwucXwpE3c7VBGyqm17K0esHVNfbvyIknPxg00iD5CTERNKtX2M9G+VYryWQx0jUD0pZCNwLvP
aL8VJpfRrWsU2F42+SLEjb9YlfdBqDeAOd+md5x4BjwKZ04tgTU2YOUo+0ewWgkL2VpmR6+zRw0p
vnSHmiPx0lykWewmzkC+AkzRhJWmykus0r5B5KQ36U50YP0+HynO+X1vDr1HGsWOe/tVI3PwcjqV
RJT/9jc96trrx8zZQT/6bomD+mI4hkifwh2TibM2IeesTGbmctYJui2R6DqWac1n00GsMd3LwoDX
4PyAm23yk85t8dcTZPr6qPkOqAA7XaPMRuH8iTe7nGFNHhHTs21Q4JuyD5d+BDTwT+vsB3zLyltv
dik1frl+ZKazhMxHK8+apmzsMLAw4uMOkJ57iudF9TOidVj3iepbxrzF9UyC3LJM4CiLN+3i1zqD
axIpwgaJ+WrLqjTh+pqjnTEzJKTLW+I9uOwerqROx+nL7SLa+nf/ciVNELzc4z4iN9fGHQmtE43p
x9SeXsEaOBzCTANOPB6hf75zDZAVDRAtEZi/aY9eZ8zr/FZCTqItV+Pe5if8/XGdIWmGUzXP68ID
hBRj4mr+pWtY8HbMx8NfQ6BGifzjtSirBeKWcUq/e8nxiduBEKOwzrPv4rXaZv0wOzV3YXnmyYBS
nzD82nSxFKOGw3IZ5zd7vUcZJ2MAXD6uB373UvktDZc0kzhn88ARvD8A4cf5SGTA3UeGQ3lw6rmV
9PygTXGe0bBGf/yXvFYjqo5ILxPVBJU3tOdK45uIr25eAKenkEugjSIvCHBl0zT8e1iDhUgVDemP
MGjS6Dm4A9JXT/S8cHgUIXS+8Rb//yiWM3qf9qibWOXusQonuCWfnpsnR5IJxff4P9zcWbktW7YD
9JEP4iZSlPybaq0LSJLG7sJ4eSX/3fsk1hUb4CFdeDj5DnNeZEQyKT6tRVgsJmggSSwTW5mI4Xst
LGaBp1lgk3eSTyWJTx9iCeRY4prc5AlT0eEg/QX5ODHMxaf0fx5Ss1QuvJilhCdYP5faWjk5Zjas
GF8G72LCien0ZOKCAkJwAX9MCcyoyp08zvFyjrUFyW0jld4myxF2LtHEzqJK5QGs3uIdbmwegMgL
2UqW8Th43NVtgs2SdT8FSJ481T/2mQX+W2+JwRp7PcJpyuIt1yP+auFM1kd/RUrbMbPNZC6Zqt6N
/SeaalXyANcmgSlLUZX39AizUzFMuYSpOiKfVnPeUAcdgpzypk/gUxqjDq+Z8YpDlUtBX6mm+1BE
rw7BRuELXWGE+5Tw6DfIL75NkaHacQaNVzVvCK8QVaiNJUgf9/4JrZxdNCE7csyIj12V+JE/CW+T
/dgjeMPSUSsdcng2WO8FvvR8UclF/ROks9BjH2b5zBu4G682t3invdELB/lzhWzGgUSksRWSbpu+
AHMG7ZCnzsw/P5GRQNtApsZ7FlhmmeYIUqlCodbB/0/z5K1DDCUVpBFlsC2s3WPVNlitOjKGPFFR
ijT2TKJlRrvrvfcnjX5XveBFldFBMROZ6PwlLOAxNGSMsOxUyabUcF0qGDM8M5cFlndcdT+zMbYs
T0gAcB+TTuF0r9/C1VfeoWtlDvT58wk4Xl0XV+GerXo7SjfaW0Y6roipVn+nZ9QYtbUuPsyOlMOd
w7AWnf/ZTkgMP0O84Az5UkAeyvdN2RDeEPzM3FgANg/pRQUO66gq2hejWht2Ei7oXxFjpibYCh7l
2h4aeO2jqAYr4n59vISMowq/k8CWWlJXZpgafhKebq/IamCypY902vZVjUrnSqNIQtQ/mO3P9vKQ
qghyN6NvXU0/hIx/1J4Sya3IHtGhiTbcaC/QC9jBpO2uXIg2uC8LWvF0Boy7Srjaj/TMdrHu7/m4
aAmEB+HOYinH1DPnQaeW+G60meHxsqaMmDA6Qdmo4q94qKya6J1Lq6aRc553lOEQg+imv/ibWLYA
m6rVaq1yPcg3+Nfj6RFrZIoA0ShPUBZ143rlYlUQduR3L32PGQA59UPbfHKbLbiYBbxd8INTVPbN
zQAeP1ro9tSFN4aph7js67/CdoeuBJHsPXbEr2j/sQ/IWLUOp9HglBceneYrQvDvOTFvwMuMRACI
hKBFb/nVPNZUyqfJZbRzn4/mMApoT6UrMkiQ0Ff8b37znWbQjlg2dSsuMf6zoIgHLA57svUFefJG
3mLk2dgSKel2O00wY4jcbQckGCPeblfoSBUBy17xgoBiJZf2G27okBsL6xakh2CIcaNipmI8bQPR
BpKLmYDBsJUBeCbO0zil2f3cbAHfozLbBwYEt/7fGcJK7iQMGbnkehFHXRGD5V+hPzc7bQ3xKiJe
MzY0tTT5RAV+ob3UFYdCtfl+CsD83LNjUmiE8YehdtiZavVYbyXGxABNcsaK2ARuJ0ePLNxv+JHp
DhFNMJ80XQ7SZ7KWk/kdX0m4wnXu/jtn3QjAKa/0TFG1z4oWP9B+dToGDYeqE+9JZ8+LcqhczEGe
UqQ3qNaaXAiRTPj1J/6BL8UdreKlmAn4STNOoDgUoB2plyFhcALube2X0Ovy/LcYMSpniD/rxIbb
36OgR6K6DHwt1H8TUJ2+PBECIsxjqsEtOUULO/jqJ7PSBvdhooMDpLZLrjkYVAQMOt2fCqrWmG7q
92vGV9040nx8hMCbq7bJN8rE3VRS5CosgtRMrG4182nwEm0N74uxlLcypmX9Ee4C8F0fOQngJOsF
zdGCsK9guUw3syaNYs8OPrrxW+qOrFFHVmMKjX7OVr5Hp6R7ewpprw+tK5QFB4hEzdKPhik3TX2o
WGukbXiyRBtVd81udoX7KWh6aT6fDtvgaAXUlwpdmkiuOu7MQxQFsOFYqE3zNYLTom67Q4Q2ZkRY
hr4uQnLRTy3QGoqvI6jHvoai3R0A7a2ive6FzK8YeejWG5blwFeZwOurYOhqswo6a3f13+9s+sME
HrYyJ5cboYOqH/XgFom9JTrCC6ValKNJNuLso56f1DNZa0vim+cIQ3oPfBoQIPvp1ovrxsATHSSY
W6PRIXNE5mlQ4JefGGEdLG0UhfQal03GSGJzS0XyuKubsw1Ya1MvrJU6GXmGLte/947awC0uvwM3
iAJ30Dbvow62RYnTKUhZF+Pf31jPzj/LJ0SdDUeohTpXAVG+TMUVKfKn3cDq1L8SrTEBcLJyEWJC
wKDkmODPnibacTBwEZdSVwJfbhr85hLBlFAyHgf5arsd9U/DfXq5GiJXxwtOze01alRUMP0rJg/D
8ouFgCDHxYGr3P1WlYtqCjf3ntlik3JQTycmU9Epy13Hjr8aDSE77zFBF8hMV9FT5vlzu4+9m/cr
A1qbIqz0ux8TpuNvs5MueSbQBvz1Lrn1NHCa02trbhv655rs8pa1pnVnNjWl61515PkgGfRy04ET
kK0zCzJCVTQ7w6kYTFuYdNF3/kZWYCeQg7IfpAAHJCnWLBZjfY7ujDItn1o0YzJEq7aJzhwItcmf
NZHE9wBaxn8USz+4oLLGqLGf2yOdycktVRtzkA1VwRFm6ZlTcpGKEdoWUbmpa5Zdi3VDB12QdEvy
F8hnxUaQ/mbmXn0Z7Z02aKJKkiDXZaOk91WZ8oNbADhr9FLw2VSBWE/P31hd8bsRZH7G017gK9zB
3P7I/crvvOeDLCtAcC0Di/WgJ+Axt1ANB9sbk1Uw4LLBgEwst/qEJ4XSJ44R//lA50/H5WlMKjxa
2bUtBJ33c0SqJt2dewhvVNR47hsf1shqhS7uumiLxHd8qzaHcdrejX7XJa/K+nkzgqsA+1lS6hJX
I8WLASPtuhD0Dad9DcaYfecDLaE3UrHL+xUBUfUOJ9pvQtiWnrrkcDEnZQoyPX2cK4I/2w6H/VHN
RL/L5f4g6PTc5au/1FSlCTBt3lcr+Hrav3ApK7uOO66D+H4UaJi9eTwOMqCzdsc804oCd3dWCh7J
l+R17RYKBRCywMReezq5dhyL672TD5TMnPbVK5DU6Yh6pwIVFM1o2iLKcrJJboruxh18AgvWwErj
1rVV6MF7nKrr2q1MokYikgBXnKjRt1Bpntzlzvmgi0J9BL/80u+gPiHbUy8Ndyc06U4c+f6vP1hH
2X/HhbzwvczR4wDLuCsN59KLyNupY56oZTNt/iYTqqRlWIEqWO4f3BJBM4A53Oj/jfwras10RTcR
fLzA5jdfnzt7rMQStJA4rJlo5oOm8KDhryJG+M3+NmCnQgO2F7nS/peHndefVItwU/z1UX68rnrQ
kRZObuIytnXFgusN8Y2ldRVQUFtSOohfeNYsgClPQynYn0ulA/MfMXD4SY33PLRntFizejpd8Iri
TZ+FfjWnFnNhfzapr3/g5fJ+Yk9ur7pkOSSVOzRyDQmQ71g6hI4xK+QRlh7uAwqu317rBvmIX3pA
VP/R8fyLk43kCYHBCTFZw1iFZG/qDh97EEB3NE8MVnqxJw9E5sF9CSfdN+xMZZOBchuW+wEYIX4W
vl8Caxf3FGNH3CcZJlepJXqOF8P+zAc9Ri+MXy+Q3nGopxZ1LPJxwCcuU+gqXRp/jI1Iif0aZNqw
XwrvDRGOolSglAcLbFLMncm7TpLDMdrwvLdgz14GiGZ07gmy3RBk1qQJ3yuEJ9OYSs6KcFtvZMd1
f2ZWjBoEiS3sxDYwSehBufahxfQPHtAv9WNwsDs7t8VJflpwZroj+cGT6BAhdYFSD/6oxjeiGERw
0T15vZdtsmFiWONC6ZrTchKB74aXKq3evB3uoCnyrhc0WKHJ67lOkIsHCQIJnGxK3TtPeG1+6xXL
h+6ANV7Nh7Tjc5j+joVP86HJglMcRuXWXLs5sn9+mEvGQoTDUWYp4qlQP/Ojr1mwRUE1/fFw4mvy
SufzSCwbxtdfHLeMAjIX+locJPWia/ehOiPnLRWwwlk3I/0lXlppWXuwzVHIQXUGnn++/xBiV/SH
v8vdrWh6r9hQy5mMcU0WjrShEZZFZzKIbPDDYGsyegTF51VuP9ov7E8ULB0HDMvStcxUH+k5enuA
+EwpeIJZzFFcxTf/682Ouu86Gkep0JmI9wZb+ehAnB5TwXNQbqavtuqLjx1dtp9HpmhkiP3nHLaz
ckdxyLtOBlm5ThsXQcUB9kwGSCHyJwloY0VfQ1ygUIG9KHOHgvmO3CG6EybBnk9x5U/GeclMi5Qe
bgiqqLy8B2w/7YWrm3hkcIFPqhLcYvukF0IUYTL6etJDjxkrlVLUEqla2KjqcspVrxQCQbOYsouC
yyFabeZb8y1F71v78KKEPpnXeb1EL7hHNWImaNxc5WKqf/9CcKWE/YlxHeAAdmTlB+NOZZ1Te1gN
cEZbCFs6bCquSdY2EY8Yyw2Q4LkJt8JMdjOktLBCh9F6AZb35Ur9EQOlvtLPwZx2RRifVnzqcZOJ
7Nu1rX2YmvvFU/3DaLi3/QthIoTdVeJFgUE39jlWtoIDeJg8fH/R724Ss6Jhi3EDJkGI6Jn3uu2U
Okz8QETguhq0NdKp7Td6jV98kSI1zlzZeL/q/XKoykr0ka1uiSFMO1GMBkC8wHsor0UT6QspdBrn
vQCxw9u4bk0qaE55Uk84gb16bHUqoztB1w7lYkprdDskehQUfk32dN4Jb71QZswR3OxkYXOevfg/
ltesXP3oIvQn1OERUjpYmGtgyakM3EpRBjJZnWPg40xeCRNrZqxakA3HdYi8IIwlJd/HZMnEyLIA
aIVJV8JHIgfNTBjtWMhJzPWgVUvkglAefU7aEhLBg3ursAn09KEmigpbaZAXuyI58xKCgFfx6z8J
NsxV8ERXSqkMUL03q4vzPQ2e4hhVtkz1E2r8AtdEDXyyp3D6Xf4z7dzJfkM/VQLNtGCESjI1DRBr
LZNb2c0jqIF/PKTdvj53Kn4i1eVuCG5jq2hrRmwsXomnPYzXaPpi4/SyyyH0Yrm+zmfbBgh6783I
jfZtXZD0QWDlacTBftMKDHJgFYATCro9XbJVcNqRpz7Oz2UrDP22XcIPMO4ayIr5vByTUCrWeuGo
fJift8td/6BIWSTiEKfSDNNCACO0B8BpZG8HSqYSiqw7Rlr62tG6YH1KUHcmc9OIcmIpfFWjfiTS
tgEvBRczlgU53rlThaBXLHJ+ijJJCVlJqOWVtuo9B4Uvll4erJOaB/tGNxYOhdKHk2Bq0YICa5VE
jAUnHLD7fUyw0QGmp5uKYby+B0x06nhaFtxvRcqnBuRTJQoEmWs9SyNLKhHlFQTSymGUpCNR4t5Q
OUiMmrCmRQoflkzTfqUU8b3SsaVdzJ9VUs2zryS+HbHxjLCWoNoWUgglaZKbHSOVZ5v+Wiqunkvp
AInkj+8zYg34Elg99BuyuY8+QT1OSEZEsodV8FKT3PpJ/fr3znu73p6OvwRmKkp1s3TXurgXwYOY
W6V/fU9aPE+Q1+ssfyLvhRrDpLyc2WwlS6Y3lccBAYia8AK6at0J7RM8AGK+OnYKfZeX3f7WXxBC
rP0nau1VT9MT3kgdBMkdOaPTl94R0I6g/2aEUeKvnKVh6GdBTS0o6CD8PKrkob3P4VSRk1XZOQ8r
QYgic6PdTVhOWVJG7c0dPYboJ62GLYzaGvr5M1QFJCy6hrUkK/ZvsIb8B2nra78HoLtpdu5wAHO5
a94G+y6qCXPVpQVyu2rxLKnA5/d9M1sBUeVm3Fpd5s8n5br4oalTO3fdhwYfoMf7H2bt2h/88sFk
fwD92b7NruflV05HarZqdZRlmKdQ/7PNv81OZ8HpDxMHvqhcQlqTgBDPFwE5snfLm3innhcXKfB9
mpH9JqyWwB3Uu7or8fNZZ6Xm2iwogQTwcKD/2HdKm3QWsCW19g4Q2YTXcukK3lTRWerZXCapP9ri
oN+hIdFHpdZDq76kELYZxAd291OLGC+hMbDHvtmC+rOVYhNY2pmct5uWexfucwa7zJf2sMYRLseM
MKIFWZIzhw21NBx/czVJHXIL0YVvVXhNChxW4TKEU9w/eKrsjFdd9f/WoVsZ6psbGVIk39WbE8Ex
Z05nNF7P07z7rCbADNqasE7OVd/sI0yfka6EE3hIsmfgLEBXf/2FVw7a2F8KNReQqqWZPtb0b8Jm
eqx7ClkIcDn1defwFIwJdZnXrPovcjA5rsApk7ZwF2IlHYQDO19/Td3WSj4mYTX4wvqRaWjgwWiH
Yxs76tmR+JgyUtcDgUsMOMiF/TJ1LU34BBQCf80y/5zbSRBB/5oet47L0ncIz7JKUBCE1mTs9zt7
4K9M0Fhsn2Oyr5g+suKNZE5k1/xxR1ENuTqUwfsGkux/7IU24wzkd5Z1+iuj1ulshATe6VNPb0F7
aFwj/Btm5DMyuYU8wbWODzfJZM0YjrYScxuR/BK/S5auxNX5d7/x8sV+aYAYr0HCdoMrqdYiYFBU
dtT2aXx0CjlA501BGpbivDKUteB9Gt4sVDvyaLopcmHzoYa/yKOq3Yczcfx8wQIY41I0I79BNRhB
lomTrfhuHiRxiZVV64bIXxgKvg2XsocM627+23ff3nswpmLeSq6Vp08KNMt5853JZz7f82bmVuuv
E4Y+MBGSZ11eA2sL5TUr6R/BypNza0b7/JPDGhJDqtljTk3c1sTXAKPz1K4xxGkzWzNgOjdUm/HQ
zWb/vrt6yrhPckxaJCmGZF8DPif8oFbb1BVHtFwZ7CUIa5BKWAoGS6gorFINoiRjo7m5hVGt0jME
/vDTIYdRqcXL0Krz5t0wCIRulFWb+e0B+Xb7DlV89xC3NdzG7iClL9HcEqdRHxZ1I9lYptwN7a4e
QVHhSlXssL9saLwlVxdKrcogD46ZQM6PQ1dZAqemI+oPT/a5dFJdbdsKai3VZ1jNESI2n88Lp95H
mYgBjlThyz00AcJ9ozkEeWnFO96EFDLpEIlcJSpuAcnuIrFsPlaOC+RnVb003CVCAVJnEQrnGGVc
xvOMIEZRefXvWGwLR/julqQcwn+3ZIwRgIR35KNrgmIYhF+45MhTYcA4JQ4/NuJCbCI2WGAEBR2k
dQfh28Uyw2kBYiGUNDOP+7q876iJC9SNDkFDkKmx+XKMxiOvrT9z8AnfEbdKOwFf0LI7zF4jN1gG
3id/v8O2PzPzRaYA5+FSPJsL7CyCVTMwkWt1kH7PsNMXWf7BkLKAxF4cnVZERCHmarwUQIqJh3ae
FWOJ2WXHY2mR40CevIppvqpUAO+FC/TWre8hAVFxGCgrt0xa3tQgSTXDnvRdErp6HvkH/u2iQn+q
UwwBiHjq2goZs2M0n1B2pbXGGp3GF4Ko9ko9uVUYgfMySfl9pux7EDgscmC8IDQEFT03it/3btuw
QyJICTTVS3BAt3Kjzy2rVBhTKevLnb7G9AsF9vGHIn/VZAjnmUPxtbUuE6uH+xJ+QJ7Y2kcu9eDu
P94dFQRkulYusO/dgNdjumVw2u+aB/yjv6rhPAGPgLrH+z+6FMu+wrXoPhbb1/Bx9kUAzk8eICHu
tzRmHjNi07IEDsE7eJQYRClKqhqBUWMaBcBGsltpcPnWIyFg1zFTeaodTx7L5eF6G66CqJR+Pk98
pR7YgcDda4NpvZU9/XH8c1ElU1HAsmM4t5v+wg2x5lXnyhQSX8rJHho6lpdS9rR/BTb92PV92Zzx
mTfy4TMzAdrEOlLA1sGZ/Q4l9aWDqIHlGM+nvAzpVRlEiikiqBpJN/vIQZ7EoCQ9gjRIBdd0WPgn
fwqfLsTvsJw1+QLv1jEGXZjoR436ZNDUCDk+5C+Lbt0TPFR7OqIqHcuqhIfvUnBjHfgUtYsqHq4n
QmFTmAmAlJT/mb1Oz7K54c/4O6QeWx4R0PlJaSV/+U8fdtdQ61fd0yTbXOsjOzoTASIgvB6cvdhC
tUkV4wuqdddg1H2dDSeo5dvTcndnLeol+BOlzmai1IW992KewAQgBwU0ZaStykHayQX7Tna31jyL
4qNTyaNM+RvTLC/ouzTCcxt/eJdzP1/0/W3xLAXWlH9FW47Qo9+xg7bn3nkzYTkYWxqYf5T8uXbA
uMT094Hyp0TW8mfdIhBZomb8lncqeytrYHVwSehXq1WojU51s0Jlmt2AR9eowkWPXVBowK6bnPdT
uIKBhZn0jGwZVqzybm9VxYJPrboKLedVD/wNe9g03y16tM4uTcnDlaokVlYZxX1nkKtUAGDewVtY
s2xMW+iSPe7KxbgJc0FbW6F/Sk6M1pQSg8taG/mgWZqxAing0JmdVmWfLH7iXMKZB9jgNqtpY3NN
wNrxiHbkpNFhDvIqwUQtvjUD79Zg/cMGJmmCINU5llZu/mVdlDX7HPYH1aXj7nyOmA3Pltbdhffg
/fM/dxXQ83QPiDgN70ZAvUOho7PaBpqMMXHJ+S0+1b1FPwbRwbEFW+fWD1pZQxdGXy+o0qxWbggN
g4L8sOfxWB7kw9QZfWcTbjWjswqyn8piIwYwLry/B3fIxXXx8WIR8gkNXUxQ6pjbtwsAp7FDbRMD
Zyrhm8I33kleURwhE0hTHedy5dMNY4SBSDXQd933lqGAvvAntynb1Zitg8AVfxhnSwyGVIOcGQAN
cxovjAz8nWxalamnqV8It2W4oIfmcEmNLry7JtX0MeYk+I9BWiU4QuMXsiiqNJnd0uVfq2evjPVZ
sfHV+kKzEvySgUIgW9Tze7yPclOPSBFzK6QIcRcZ/5TFFZwTLBi9/jUTqv1JvdPwgJn71Q7vxpnw
aH6a1rh9jZ3tjrYWjhUNuyY+NVF3N3OZWzLDELfar2dWj4i+DTQjkC/nTTJQzlDwA4yGckIAQ8U/
F90IZ6HpdfV8916t/Oi7rRvHb7fC21YMGj0igPWCv1l9zS9w1r09x/IdnKyaY8SJd9lnwABwDEJ1
VT9VD7TMEiu1+F2inuBd2S04VLaZeUw2h4PRBcnT4dpn3kG+iJIYqc8Ce+OIxku/j3POYE16M796
UHjkyeX09sfP1XdmENT7OrB+j+t2y9bZMtyymiU/Q0so0CSChbn2UA361N6fMtE6azQlCpcQDp8U
c0LB9r3bOk91uJ3/07mOhctw7+IDVKc40mvb+RNBy8yUFIgKnfIjhxsh1+v0ilHH8+LxkbDwQEli
9oAtI0ILV+ynM7ZDNEX15PNsC5PWlX0GqfRzUKjeosvlKRL4RToUWW8zQiVT4TV3Se8Z706zV6ZN
RuNkMMObeQJ+xmVQ4vSgbO63nGvS06WNoraOAfwBWaDqX+1Bcc5k60Q0ua18BhTbhoKxMThBnHbx
SorwBodyeFrCm1u0fAxil7MQ569PBNx43ZBS2hkg332q6ZyK7q/+hYgFRmQt3SmD1l+DAHVvhYp4
/E/nRab+JntqNCdYoTj7smWrOKpkPMz89SBbrxeYnZM4XIcdBqCVUKWKT9IRId75xQQBB+XGF47D
U0g0d9YJjbOUfYFtY8+2nFBWtGN7y2U2xxJquxqCBBhLEvQqdWLEVFm91LyMB6wqjCyE7jne3RzS
2xe6xJ139jxqnnJBl5Z2fkxLmnRXqvjwqa53Ggod7ZtFOWpkGBWwAo0dHwY7x/74n904IcdCeHI0
Ru11u5kjoiixz+2CdvUJeP9T7bBYBKW1tuWvt8upQmhUOmqCt+woswBgZHyHVaNo9jgnOnJLiBJJ
Er+1ElYFECO5ytPeGSEWOwNIXcJI8cvDcPcqCoQmt03/OIRy71jfbEdv5mKBeEW/QJs0LF2OOZQY
dliPVN5N5T/yFTQkSbSKZlps8SBz0ZgGe9MyHsFv45YxFNvuXwMJweSkdPP/3L+58et30LZJZkCS
o7woXd2Tdgygb2AVp9HdydOwfryjbVEAk/Ivn+rssdT89uhS1cyjYwFSgAQtj9csoiecU50i/pWc
5N1+4nbJiHWemJzlW0tBAL+309PUmGbtoOl1sw62HkqkTpToszXKdDyBVHnySVJCmN9E5DXOo8KP
02B7Ip0t0X2+7F9kuypK4CbyVmFrSFPu6Tj55va8emQG6T1B6akaRJhi+kQhNbYJQEqFCF0ZTXmL
FrVvFsfBobQIgislc9ts8zoVoTIan3+O+VOp4j7rkaN64v5GwsecmkrZ3X3kxAhhDKWUR9ygjg/l
P4UUh4/yIASKpZNactmJy/M9j1NDGj9vB/MeY19A7aomepyX1L7s0O3CYCuor1RAsUt5hCczXCNp
Y+RXm3VcLQ217pPfZMo8h4WCOmFtjdzMJ487/3EyAixsV5frdHh0ZqXm74dVaLW220Xv/ZgNbriB
IY6QBH8rIdI9B+DzoQ/xhSHpEAETeRLjhzm9i3q0bZ+9tOWyq6nRjffqmtvLU/QnPkGB9Ej2OziS
xW881xcwWJKSP6uGbv8eGop4ulx3LGlzHTnRDYsTTVKXpr0z9j04BdZPCXD7VYxNz7/0Cpzmg3AI
LCfvJjXWJ1hxCQpPSWhaiijRbnR3DgWinLNyP5fZPCIpWtB51dHywWLjFBDsIfMKWU6j5wBuMgv9
qI+aTXthwlNocCa3IPBONIm/0WGtXdIHjPJ/3yDqvkwWxpP+oeY8YPAR5OsBVnmU+LgyMLE1/XwJ
uA153NBtyoLluhI3w+/BF6uUPLz6jsFdp7wb/L3VVSeQy0wLrZuRAXO3FBXptaJ2k8Po3zpIdu/y
9xmgg6+cpVUTxVPN/EAQvYxwkmCNuT5+lnYlFwHONAWunIOk6CGrjPE0ULhDBjDg1EcMKCWweBPn
ccBXEACMmWsfSa0L6MyHWKb74cFpkX9HOSO3nfaJ+AfCwjJXdrZF18sKLqUl8bJkruu1inFCdC5f
cWSE90/JbcdtIhOfN3wERjiDSqoINNoghqnxDB9cpTDC60BtkcZlw9SRnHIMvjIy1/+vrsYXDjUi
3hiK/Cu+pZIdOguWMs9/LdYnqVVakGBvfcf8e72r0Pmq2KLHUHyHV4p2phl6XI2WCVbCkoL4nBoC
1v70f8j46FfvgFwQuI1pI3oKrp2+bPbfGQ9LCiusCN22TOnkMWGSrFlSA5DuI6PIWqwZGlG9V/61
dehyOua7e31shi/zaQOnxSMjr7B4/d0fAGC408xS+Bt3v05z2/KmWyDOmLiO2z0+p5RFOblkFb8v
7+8Q4VCDmOwcUSnHo7Zit4r9rQFHecJeXMRWPfWzvw5wlAWhARjrXek5uTakV6b1DIsrgQuFBlTC
sxNzPEGDiildZQzIEzsy2XxmmsR/8EouyB+2Dg/xFPNBrE3IK+es7ZMhki0HS6yqC4p9KftDq4bu
R55OUcgjOg5a4WeecJOWxzMoYLijngMuC2cW64aTPivDobEM3bLV/MT5x62eRPfQPzI0Tjj54ByN
okUyx0whbiWkysAckdjelEpVeGOwgzAS7kkR9bqpPMep3TW1kdq+V4a/vuqc08wZgDUDmQQ5j/FH
d8j0P69TV8XI7hZkqftFTXBel/uW4jzJfbOa/kqnUeQMmpHD+s0mqnQRgE92q2RAOKSNfxMoYRWX
INQe0PWIdOon/ihtS9r1YN42S+RwQrJj11PG1b4QDbpWnpZpWY9OXOLrmP/iizeZDj6F1VqlknfU
69rKj+x5F+XdJj7hGkmRYAVladz6uW/Sr7GYFuao1yi6fB7fOdcgx12w5Vousz1T+6SFTfT1XSxx
9LC6gbzyP0tEga3tEjm7ZhY5kkJ5D/o/j6Ha3rbrsDLlTLKMrOv+WUv0zGVEt9rvS8SBiWGa/f2I
fAiCL864xnyPiiZ6ptAPcEWYfuW9jffor41O1CXKdz4gs7JvemECF+SgDqDowPZb2Q8FIqfnm8+a
csXnfEMNEAqVnYES3VWQIrsFI81TzvYjF+POazL0xyfEyagPPaCEMh/7kBWXh5tLFZbjGKqlUmGD
rgUuCjXEO1Bypy23Rl29bZ83iYjPd4p62OaMgUtjWr2n7uHQFWGlTKFyuByyRVOwBj+6yeOP0E0V
4Pk6D4oUbkIxsUUN3Q9fTrS+6ArRQG/6l/wtl8jXmgLCVV3mtJWJzhOEUI8HeEvdd2LHgs5a8Rll
8C20ortW+9d4V34MEo8faNLeV7UhObI3SeLaY5MDAlI9UJdd/0Xoe1jfsi5Pl1YdpHi4qMuHYYR2
3iqPgaZ5tMZkcv/by+zv22WpHlm4jSfSil6ts4uazgZuPZw9emO8TmP8NPlmD7UEVRfr4vT/Ur8x
1Xw4S3uLtzqTWtBcsOBDRtJYpZCjoLTTswaGvasNzHU7uNbMcpnC747BSKzEBa2yFd58G1pYH8s8
vmtE7nrZY04MIBtRPJoxVdLAnGk7qi+SPmd48rqAwtmWaYQm+TwYVgBm/mjvXcuKTmkDpVyKC1Zr
zAQf03t561tbfRDAeaAmXO8a5anzCnt/ywxtWiVeWflr6H0L7OLMPBD+VEWYtuo5YW0BqGW2nC68
qb6Ni/QiLZPYidfLlIbfts/i/86FT0rSpcHsEh4nZ64LK4IEQnASSIKebsMkE5O1Ssj+dWQ2mXxK
59TXMAG3S+iq1qPoX8VBosc7nblIsmJ8y/3RRmNMTXJ5n3muM/BMIXYpR6oLEKtvJ0HZ/iI8GTk9
iCSBrGsYPF6YuY8e6lS7NGXLL1qr3ZAHD/DHLje/hzHjYZbNV1Qnu6CU8xu4d45hZLUKBpCF4zeg
xXVXF9/w4M8fMLXuBUduZQ5HVkhZHaGXQ6dXwIuhzqFnFcuWNSRo8/Qt+n0dnN2knhqPCq4W1HmQ
tFK01F468ZYW+jaXLonCRnSQNIUo0KEwSRALA6M+6gt3AG995BZRQn+LeIqG8lm8+MK8DKCJ2Aqd
0UjnuLNSCo/AWASRENdGA8ytUs/6VJzdrgZ/4AiTkzN/pJY428W5feZubvAaRlAVLQxUsLIsdd3O
TJ1kSHWaxBPzM4zgSu/7DWAB4QsSn0fhCIkg7TToqRD9fjRzv9QUDFddS81Pk0aTOq0zeAd/B8OM
fTAH4f9iqjbHbxHHZx/vLgOCEJ1BQGKfKRVnpNYbFw1tDRZqskgp1yZXzBpmHhivV9ngZnFLQ8+S
labbAAh/k6ExOXV4C0sXmHeZx+zO2nJZFWvwwq4IhAsWbUuezcr0Kq9JsPwb6wbvigw9mJQd54+d
DHeOLCUku3KQnalWbwoo4hMsh65R7MGf1vHetWo3o0Xa6mJ2C0NINWr+hMiGzv6h2uoy5gF39FYP
czPcLLKOobvkKp2xOrwB/HZPvxsrzdhD+HtlRpOIf6JCMYRztWnuQfEgPeQSNHZBYK2Y2zkY+U9x
RJZaWPCJVjnwhYfLXo67LUfTum3gh7QJ54BRrh3LH7lRfBxWCVyNpRVUFjHNyz78rqRQgsJ8Ri9i
/S+FnD8R5nMJbgEi2R2bR/mmrMMkiSkxJ3Vd6R2m4XDMUwjvBfbSmOp5Gs8R/naD+6o/LN/C6kIe
MEFspOsW/dCZ/3wwUFvUgHWDUYrMbNx8+lWnKHeGS2f2y+DxcVPVA8a5swbcvjbF6ZaGYedvPX9t
CDd2cSxPS149zmXdVUM1ZzYx4Z0aX0WpcVl7XeRdP1XF4/mnQ2VXcspOTo0s+FVWnND9En5maf+n
4hwTb+iS+EIPTPS3q1ggTYc3oLCBwJtQrgFfMa8b15vDgp4l9yQpVKw0wwBRyczMWAD8ShNQOGXb
KWaivAo3uncYb6F9HgckVEHNB3vhEgPQmuuVOmWGwI5IGW5GCaU0mNh2L4bmdoJAh0rsqFCb5All
PB0tPP0s/nEktdtWnHdkVtQbLGysPs445NdgXBWtnh+85RlP38D9SyoPP8LB+By+LxUWLKnCmXUQ
R7QTO/zp3YhmoeeT1+oKHMHClRewtqZaMvghJxS6fKSHDfOQ8ujrqf7OIVRLtaxMVkiIpHBzXdyf
PYKz3V8komlQgrdS+SdfGG2tLRMk/RgLH3mYUWJn3G4rfZm5BAKFVV1Ugj51WNBV9i2NEq4/ocCl
D2c23L49e0bM5J5OKPGHOFyhCjAM4K/BUTDzrXdLTwKrz3B8hazj1EU0/gq96ZYB2/OoMaQG328b
IqvjPIkv8qM9gNA95K2d2+StiVsiUx7/FzNtGYS1TvkE/Rgd9lq0TeFMv/vxPeTPOhaPIT+0DL+M
zUPM5MMIeRMf6glghGBHag4TfEKN9FOq9VQQZcyKGnKIRlJudjEOgIvjbY8F32jaaqmQ2cIjcL8O
aDAaFuhxiwd04k93C4XbwAl+H/28ad0ch/6z40aNT3SMYO+f9r8sGwuiI0HHY1Y91vM0X4Oh//by
Qw2p4bdeG80WF/axkLFNLg1mcK6rcOyAsBi7J3Xgh6Q7vPNPyJ+Ybj23CW3fK1M3we2f6mK+ScCP
74wmpl12QLF8RJbgXj673RIbhI+cczVGjYMvYtWVrRjBlenX9krQ77XubApDM3uSmsLlx89xXFU5
AEClrJjKAV0s+3zjHrAh6C3zFUIDGV28jM8tuV3gisLamd3qcrMyMNPr8P8P0/Qhcx+91F/g+Rau
+wvpCMR2vtHiFRBbzZ9Vjvscc06KnjsTXO3p3J5OCSY8Z7T7DaafJTiOOHAm+3pCp4Xwu44CxcsB
CKrJQwNJVS/vIxI57JuQdsYfTkRT+QtSk1G2RtH4AIwmoqW2B5ZvwncgJgvaILk50khtvUJeXHMI
yM3oabfSYhnaF/m5kYlezv8kBo/pVcDLH7aq7k86MpztxZURrWdf8aSSJd2DoFIROYMifU3a0n5x
OeEqVojBo/bG2OqhE7U/1+I3XU9gtc0N5Iin3ymwhsX1jURS013QaAzRPM5/eo4WtQxZtKYzobVZ
X2oEVrB+kByFf25aIYqYF2sWwrf+/2SOy69tiFuj3HTU8hsV22DEen1NvCnEWEDQBC54a0fZTgSy
qy08qRw1PFHJcVAfwAX8X8XiW959EpAaOVWJWxX/KElaoE4zC7Yob8Yb1G9yguIOJ6ryyutMJ/eV
7gjbPBISCiI75bqQRtlvqWBbmGbq3IQ3PDnaJA4hjGP7NGzCNJcj1hU0Kr762ty3fqbXoqo7q3Io
v6901g2eAVk0O46KLcXhsBaWAWd92wR6z8URxieQz5aWWMUDqqY7nzE23oSZx5I9nCMaXTmpEzNM
BrBDU5CfcJpxeXwRIbQN1Rs5QYVracUWvRzWi5QC1h50T/tsNX8jLiuXY5F7RH/ZV2L33LAYRcwo
fOd1rBRKRDqo2T/YahhxZiD1a1kmotGTx1/CJXY3mWlUnKXyckzcRALzzrI9QlilJZS2QAqBzjnd
TIubIl1B8+B+wUProuqcSbFKGamSkMYnFCahTGD/0SuiUmPK0xD7QDpm5w2m4yGAcaEfphFnvu8K
TEJIwBOZFa7iz/myr60BugScytIttRW6KXf7eAUrXgAuMgDlMz/LodZZByDiIWQcxfpu0zFSZTqy
u++gN3ACCEt1svlXRkZ0Di+QI03LmOw/ofOk5iuwiZ0/qEWFHqb2vAVtbBaU/JlnKH4Im9IM1lph
GwqLSd8KAHpu33hZrHsT1TVp33+WstaoZjEa6Cbwn+FcSYRz/R0YVRdU1ObBdf1RVB8T3ZtfChmL
qRO6VsJo8tOUV3//QKPpxEMdZKDHSBHLLXPnRLpSmXwhR+cNBJXK6P9PPJwlOXAAgvI02xLnaX5T
7qfsQIvEu0Hpo9zxhOl3fdPFovI+iHeYN+QMj4+OY7opXza9OCq4uKDaaoJPcuQjaOvjZ0DYRAFK
oCCokmlF/eqFsxT1CT5ERJClJ/DlawX0R4UC38cgZz0onipXwoEh+XoFkKfhNLZlizMb6tgSwuEe
IGsQyFuQ9x++QcUkFNwBJ9DfbO/fayEJseUo1jweGoBEhKrpsqkdgo1aXYlibZqBM6zZhPP+ZA8P
qONQHy3wb8YYkHtB2zY3IYLT7igxcoXwYDKaAZpdQhFXO2gd1w1QbSmRTfZMzi+KXUJyf1f9JhT1
Z7ruSMqh4V6IGB90QBKWshXsg1Otn5zDi/fAUKKNXAeomLt67hnc6mYUTVBH6lsLMij6S0eWM4Bh
ki3q9T3o41dye5J0XP0X2VYbr3WxpG0INF2UQ7e38ybYsrdL2TKEyDXaGd5xEKqrkUIo6n5C95TH
qZaDflsvY0ZQ//jI+KeeZxZDchOAM3OzfK42rwy+KbIjR6H/08rtpeuPHQN3+t6m7RwY4glMpFFe
4qlryOVZwPwK0gvDbuqukshCzNB9JI71IeX+8nGVdB0Shjm5ULW+JMCoWTZWDg5JiqhW7hdYqp2G
Ia3Ta/plmnhUt/7qJxuj621O0hbLovBLHFvqwuZHTJVOlNWj1HvQjD/txoi2LUvaml1tGprtinzK
0VVtj2SraCe6ixJ5qAQ15ywKFd3WhnKrrnrBsQ9uRxv8lxI0xXKlqZtuCt8j9hmiGUQLi37HmYLX
Hs8FuEENNUOKqtJm3iBJ/kC9NGhNRXTyu5Yv0+70yau2U90UjwYbcpTO5hiX3ZnLDPH6y3xY4SVk
D4hbP2kvaBBL+TPhttRmaEjNP2PiVzBZgk6A1vxjSksg7YPGcv24nXcHSse2t7DJLSFYLs5h5ddI
aKrK2b6JSU2Jyu6t83o8mo8OIynPlKbVAk/Dl4hxE4Wd5B2E5gHFDnm/Y+nAgGkZgGgw7wH9Z9EO
n+g/vVM/Pjad1au0HG316l8TIvuZ8/aUALmQxmYNqC2jq2+8cibE23RGrekDbQwwEykJsFFaODyV
Po1MMCvP3OP4s3Imf0+Ju1s8krHuqeP6mp8LKF0vQHfJjIP1Em31yj7u31TQ89egYgRikhVWOYQa
xAtaKxmYMNwZqaur3Kceo9GL5vm1tTYxR50/EvgqmSfYItAlfbS0kBAe9hl8FP87RGLclundA4RD
eFfD/AO/W0upnZOM/OQVnzutXzs4/EGyNGesIVTQ6eac1diInYICBSZgivwCgXbyLZsM/Jsl38aG
BHPKL4mW0xtCbCaisgDghTwoyO0vkm0xMKbVkXnLD1W8YViZJy4r0KxnGhkRms0nay1afAZf2UFk
ZhOtS+9Pxmfltb/Df6bU1i0qUuY+uHvViXmjCa/GsMR6SaGR4z39Mb+U+wEL9GYlFuZpZ/73ZDr9
kpvkBYPfIdnz8RYW4/M47mN9Lb8AeNes+1eixhl7028W/1fY2GFvKZ9hA58drgwB5C9qu1mpXBol
pUq6g3+AzSgEJ888yXGUPl8/xpPgPrX0dDAAct6kjwcWzMwnOxMyknWDpM+Wt+WfPHbY/B/9WGUs
4BXEf4Ife2TbObLVGasLowD54dRMZpF/Vh2XQP4U7Jw8jmXJKMQkY8CsyQZKSY8uO4NO6r7f89Jy
pgDp8mePu3GWdSfSdUWInkfavP+mH2xE5No4WXGAzqicCLSS7YfcOJl3Reu8j7M6RlV2AYI2cqoz
+LRHPQKfHTc2haf51ef8VikTdQKpzPup4RFWqQYg4wFuVR08d+LrbonRCVrk+tvG6kylNSIovSHC
ceGk8InWdrWLeoCtLPYV8vL1Y9mOy1H2yDqsUP7N2TUpVb7nw++mvfHK/Lj4+7gtnkNOCRXaN7kQ
XB876NWTRkcwOkwTNniGFJ0aKXmb7QYm8rZ9Z9WVUTZsaRekCLz/5MxaBeLN8vQdqV8YZsgzyjl2
oyxMS1iLiLpQnZt3OLP2Ds+BnqOxhpPStE9J/0SLLKynZi14monyCiRXdJbU2tjqH4CIaPZlTHI6
WP611dkC5p6yB3LF2XSuX80/NEaHtQR9yiQs6FWnmT9Je9tKZs+YxE931dWshsUBh0mEcM8G9/Sb
oRqOd3xqmbm5ry0TMxjWNjpkPjS+r+uZy0YN+pxEEtGUoA/kgKWCHmuhy1zxw0EMc3sLgGY+CTB+
9J25i27bVXYGB78qsio3HUEv7w/j3tAdNupjYNcpQ0M5IA0AqPGJV5XY+M4Za3TsrAJrA8+dVTy4
Ht19YtG6O8M1GTxLEzWANKknrsTcYE93k+ahGVY3+Z4zT6YoWCyf/FYrhsH9ZOOpoanoLcOomiJK
SYQ/NYYNyKCnkbHjW+9kZZqw/iFK7o3+C8fuYE91K71ReDudLxhcSB0ZyNYYqoqRIIi/ZnWxrGmW
pU9nDqwVhoVGBndbk04FydC81Q5EsPHr/lZliJKD0bLZh+80VrSWO2bX6dBN1hac/J/HZu/NyI44
SvIWSlvSzqmcMa1VoJ5V9c7ytj69t1Sy14iywOGHKeuCnJKA4YSMhXrj9n2YtiRMNlBjQ6G7qkpa
hcs6RGl/m2pG5StT3KvhdzKECK6dEJPptJE7IGXuxaitFO2PGBZFQuqzNHrH40RSyURVl4TpBL2r
3AMCWIMVKuXBMFop161Xz2sLzF7M5aMzOpohLpVT6GAjMCZT3OUiSHPRLdqU6yy9MxqA9OBuu3vC
gbe+DBUXu509HRCXu2ofMHAA71g6GXl9bnWITVUqDAJK+wXETj9e49XPuiBCNuiJdHh44h486i7R
cgu/6JDw89CoUF3as9/UcFCIWFzmSTp889IKqOBWSQPMSJcK0HMAD+ESeyyNiDndRaAEk2Y77FCi
R0xBQcJHs9x/QbklOrw/n3156UpAjIRPR16dJ2/uB3nfeu/INveHavv21WsVPauEIqd0IrRM/MJ7
yXIDbc/aBU4ns2HG8PTci6+G5uIWDZH9wV1ObcVku2j0u3HMlh5B1+/hE4SLRXOyokgELADlAZqy
/VzGm/Mc08Xgrg4z1/3CH7d1+Rsx9S4VAOJx6zjl+yWuXOwCuSlNxcISrEJogT4JZvnoOJKIDyKZ
m6l+n1pJosKqO4P9GX5hhOyFap+D3We2BSJsN8BFq7x6iOkSxD/SjTioCmMPNU8cvVUDoJeACQQo
Gw35JDBkAvS80gvhUykkoXf73xzrI9XV4yo+AxslBc/B0Dqs0T+89HPrTB6K4SF+1snGrBeIH/UV
BtQgjpEMmpxacFJATcfjkXxu3tD92gz8RYaacwA80/lq/S5cs7XcSm1BqAWSHlB1wdfLelO2TFJO
oqsb8jdll1FKRkODHLv45KXIL37jt6S5xD0WfG9MtagRD4CsPl5Eaht3yJ8o1U4roj/sWNgOpWBK
k667jzloKw9FVpGkeAoD4bI4sTmBBCSrBXPfGbzBOvMPTIU9u/Phi6PacxhZ9Fk285guD5gS8IAq
13JjWEgEgrj1OyqT5ZZdmtfyAH94EB/erWKh+YOjnDNZeDn9sSZOguNMTy0R7D/28+K58luYeSOD
8Jt94hnkhFoYVkjxJ9Ul+Bstbc4vnZdwQxmbgtLLju3X8e2CgUEd/Eam/D4N7KX0ZTXCzOaKL9bC
PaKb0MMf6h5xzkxMmDeK5E28pLKAvgmstVcWvnmVYVAWuIp7zNqzqIxiAsVdxbAkjER0y9tCN88g
drqF9y4fRsfSVND9NY9W3LR859OCxU85nWef1b4WUpAp/6LxhBoifZ/jSaVXHMhH+PdPNcVptKEa
1387Oh47GMRo7WwC0A1OY8f+WUcXV9pT8Pyx3DCcHUOZ+nHIkD6AoQKwTA/m76WRqZnPijKivz1M
7hdpALn9PfHBRPpnHwKv6PpH6PPG32vw9fdEwtrw38sTk6qLn1ZDq0ZnGTidi76EzD+EeaYJ3a87
1eI1O7EpBOBPyJgIDvglSYDB1ph844R4l9ux82YXyFfRqvQRl+sc2iHG0ZxTvkElWRyvuaIL2wNC
BDIX+cSINgyTMfsCdcbBf/rIxEDldTfgfU2eSbowsFvvZzrX9Nq4q5bw4hNYi43bOoyzCUjZrZzV
5oBypsg0ibEbvNn3+5b04pc+Vb05CvokmkWGh8plA4zgNSKbBNUe9DfvxJdkLyPl1kAOQxroT368
NyZe2WpHbiSxal5KDydhtVprlDJACttVyf3p0Opsryz9vxJXhYMlyPAo/A4P0snaICqEjoBPJwzN
f3Lhe0wYHbkx51tAREWFvrDxjHcTpRDIjPzipcrpsYiU1HD/WVrbrNHHyi6BstIu4v2CJZ0bWbjl
AOTbcC9AM8FRcaZAPwLsfw4upUOI/rEAClCYPwuvxgLvH9O6CmVzyWT8VuZ2on6ZIHO8/G3HWBMl
qnIEink7yAyDxeA7hU/yad1Nr1GVsfAd5Ka5h5TrL9+8UcR21lQoDA5jFL6cx36klUySurLMJBZ6
s/HTIUYgwg1ENEoDAToxZoxdptGlkspjZ5JBNxr0ZxZTARDzA1iT1XpqhUtJrx33GQLVvLTIot7/
Gp5r8Nvv63nLOTeqiIVlntJwx/JPzjELXLGD5vGPC//j+J80zePCj+u6Jqw75O2kJGq3mH/HXZJ/
QNwqfomObAfUL9edOHqfi0/wcq9Nugeqzkl2RnVV3rtXbvA1Xi9sgs7/QTEDRkXSuL+LGrOpHFdd
ApmTwnkG62MHjHJ5hzgaWy5cMF2ZCA5sFzT3diSs2x/KMhKoSg9pVjl0EHovjMKD8Kgpnxuj8aw8
LDwo+wdPM9jqBm7QHnWEwYFq9R3nZdPs3Xal8Fzw48vMmST79ddzueok69f6b8kF3hillUGpSTVa
16SfOhaYwY7OucjiXyT+EywYgDPY9DOXgiO4SaLNwgpTx++f6LhiFHGj5YRbWhArHcwmXdBYmQDc
d+1LEko6YnTjuOG1YcXOIlRjUHCoZyeJjZvKb+9/LsBbHL4UY3DA5oxtPr9EepGffOX9XwzoPE/g
9iXFD2qdeHGEEx8rQ0a3Ntv9Bk74Bvd2SBiL+8aMuddBAWy2rEe4vQWI9h/NEzblYZyN1N2DZREo
SwdQSjfSupkv6U1E6wvhqE+YIGmoesw2eHfJ8TbvaZWSVJ9T6580BNRKwyVvYdEINGyBJDW94eOZ
G1EA/g6OqQWJtE7CE4t7jIG8an7XWIctlut3RtBHcx/oNmIwxv3m6Zvp9mblb8oNOi0aBsa6XH9t
qkFJEJ//dAVpgxs3+FiuRClpDALkm0r6QOQuwJD7/HW8nKTXBBtodNSU2M6Y1VrvHAY7wzb4kA+c
xNyCr/Xo+TeCqDAtGU5QcrEd6cRDlSJ3BNAPodjGQAAmmUdkdhfMP1TsRvfCMQEOK22MgkDLIej/
iiWD2O1J0BntfdrtMkf/YPCDYrQWBJK6336VnHt7hcKVIYhjeAmu1vwe4H+FMoVtkp8R04cEuwd1
yZSWrFrOAF456DNpA6Fs2T53TLtmUinGThHQuxz9MbF7whla4J+VFpXt8m9LKtF4TOtLLSexZcoh
JevWUHB82+ZLQjPnwiPXCv59f4lOmU8RSejNuqnJGrALca0QQN589Lb8or671ZsFReF13vmRHFJh
GmE2jbuiS+ZLP4jwNqh27OhJTtlVdRWR5oMySv2BN5VJcSQmANSgOPPAmo0qlgREzM6Yxj8+fmy8
0l78tcmwqJR6pYmwi2u/sIvEvvf9gtiis7WmEZ3ELvZ6Jj7J8sb8XAcOySMOOMl4guSb+DWx/kDa
xCAK18/Zi6bI+RcyObjz9emsVqld4ga7rDq4+QaG4XxunymUjJFRCSGDrSCwBAtiqDX2yivG4Nrp
WOEyhFLuB7h3bEOdZixW6YA6MvZZU8EJzqIUmpotT8DG741WtkNZi7mtyIvNmyJ3HxvDevS/8WQn
O9WhNOTx1PgySPNaVHS3+KoiKTeR/i5AEbuuXJdqQv6T5XITAs2XtHj13OK4hCZ3fF40f9S1JtTl
cpVPPzapGqVW5fivWBDoAaAtJnDaHqA8Sd0vMVj5I0UDC1uxbQEuzOcOaim0qiTZuuQSdU6PGoCk
vjII3J/CwjW7mq0ldUM0g83QcNqSis5y7oIBOLmc3bv6E4XUK1s+ySy+fAV+P9JOG88QlsadJRH9
bJ7sEdwDmNoVzbWQshOzLB5AHrduFEEEaZVIHqELCvH8/fY/KspYogRVzxO5KRzr7eHm3AFVTm5q
SmYL79uXkoQR7mXD1+5itaOW6REQ89Gsv6sL/CF8U3IboWoSvnVjfZ6KHmTBH37o4QyguEMshYKv
bgN2khGmI7zq61N/mWgu7GYZTuy9L3y2wiwoym3HUYu08BnocS2nebDjyveJPdRgXKmEooynm61M
ziER9AQHHOJcORlzSF4wqVqZey4DkwpIjT1qGdA2qUhCos+aXUAq4aGK8bLEjSD1rLML+SXJ5W34
3QXnzknFx3MV7SVNKwiTiQAhfgUHpE7KmgMNYpGTjSqwL6wB4DnQNHRGyHjyCoVsm1QlRqX+4Rnk
HGjrqqTh9xPM6O6kzK/FwANm8uI9FV3gISS6WLGqHtrzVFLOfltKSXuctBRYsqHjpqfpV9b0ohrW
dAELkRUO69aJprVOqDv0N+XBe3UFoBA21aH0bwKucG9442N3Sa8x2PiqCr5ZL7T3tW+GmqplI+1C
8kxDoX65kFKh5JaevSMyi/Hg7UfC+JYkc2HnLv6N8w2YoS/qe4oekO9y0u/ESY491KApmS7WyHZF
qffaCZiE64mDjK6fS/SyyvnhlO/ncqJh8LBZVUPszYN5P4M+DhrF1TMlDUKjbbtX3wF8iSPRAEb1
LM808SyK379/43ZHFOV7IoZyPZ+OQsA/aFddXtM9BuEfraqywS7h5L9QOnRxOvJZnt7YxH1j2Eaa
j9RGlYI/dtRTg3XJhkhDmMJ++JXuk/fmvieWW/exW66Q5LFRgtBD8dfDcsGrMpmNeTYdm7vZHSiM
Tvs7XxFk5r2PwdKttq1N7h1+OQ/xN9lvFlGz3tFn4gaRHMKeVpvVbhtEHIugNBrUGaFJpUj4uOJP
QkzPvJHnWr+nMP9IIfawuWQ2FZWLtEPPdqWMh4QCVVoo3dFkMIS/k+QRGlyzzNjL414bR97OIx9v
f4fUMw7HAYY5Fwnv4Kud/Meq8mRNoFcBwFcYk5Dk1mrsi9wAe4+mFGJpjYFknnpV/bGKqQDGSbxs
QYs9WWKgloOXbSzcivxkxjkVds8m73rcM7GKtRTl/32kd689MZF++roAT2llCFvur4L7OM0dlUPv
jtW5R43/B8fV3lz/uuVt9kehgeUyObAnfDMReiShTIyFat/eOyvrWddTt+TjFFUP+wrz5WGbz37B
lJA5eldgxl6KfizXjpc1GWEr3O6GgC1NAP2EpfdNVrB2VIiPLHGBjsooIW4c96yAtIcGxYZ1oxhG
pLDe2/WV3DCiq+XJy8vVenqZ6RKICP40Gex0IWYBjnmS2QJhh2HucZNGIIYBimPBNSq3TikhUUFo
+lx4pfqumMVKHElXmZWf45IFzVDLN95JvJBdlCKenmJ0JJSw/54iHj7VpeB6MQ16TerYVfY/c/Dy
w+gaphhkCy0Sa5yoxrcTje6j6IX6X1FK2dYK8BfBG0wkgfHuvtddIWM1W1zKY0I82tfvD4Bm1kcP
CoSoi7RIEIb1+y91tdETVIhomeVfbo1mM7sEjBcPrw6aIa45ele2764jhCJ96qPLvNJ+rbqmk9c8
o6vEtJ+dQGGHUUrriUoVpVyO71SgZgkAj7qGi/LvBEhYmbuAegUytdAckYXryoYS+JgusnFbCq4X
YGLorgZfM9tmMnNZsq+VO1+lkgw0JKqPnrgBByZgPswzxD9LbN3HVvQv3Lz+cRR25Mh2oPZfnXTX
3Ybc9tM4NBiIFcrahgfunOHYPE2H0YojVj9SfNa9dd73p/30naLqWqAQMtkSG/L7Yv2F3kGi3HMc
AKfNH55UZlyTKVNxPc5EGuamfOWSEE0JgDK9UbHAuseD4oOK2dncj366a8wdMWwkPS7xTYEUQd8b
nB7QdsOBo6ZD0izPJB6wMvEa3PBJa6r52ma3fKHycx7RscewlTAmVhQf+dXd0n5ax5rVGT0959QC
6UVEA22Qbc0mh6pd0rdC23BpeJhu8jkZbb//eIgo3g7zNoJhHjSva2I96OCsHNV9vLtWeZAuKkxN
k97e2+8rnrx+exAkwLn6QwlFMRjow2sRjLb7gYmnu0bNmFSEQ7tnIZbINbq/Bs01OVeMt96X0jVH
uGGZ+NWbAfOBJwyPuqT782KoRJqnCh4n2ICkFakj58QBobj3rxn+ohSkCuE0Gx3lcXME+A7zARM2
89ibOYPol7JD447u3QaTaPUMtoGg0RtCXb0XSq6Aq5ydukTMBuO5AdoG9+nlQkXa3kCwSZiq6Mx8
kHFdcuLfm7kgGE4Jn5q/HRPHBJCYGzPXx+e+vPdrnpyakKO1wuKzBatD6zKRFFwVE/SqiGVy6Mxy
xbDTFK/iox5iH8Y56xfMVwI13H3t0P0ruhIxzHT14k8O/pxSSIMM8R5LcUIS3vz8Ar20o7aVU1xv
yrO3ln/CBCjF0YpQ/kfAavy5kj2YpsUyLt7qANnlckOcTl7zbQHXvUgqk3Uiwe5vSMD67Wa08dNK
1qpqwzsOtddZ0nmc46VOJohEdb6p5di15JkuNpNEE2BS429+s9PDnVloYvZrmUTxtZUyRgTCiPj2
ByaPNbbfkaDpZaEFN7Vp0SrixlpIQqb7+rrMDpM2ds4Xiur2EUFeBs3nZnL+ndGOGoZCAHXpPbh5
UcLntElUUtdvcMDfoAsMjuhh5v/uBGtUAd0ZE8kRBy269wGyLMDz9O73katcWsY2FJK6N/6smfsC
LoeDIxkHDBXxP878GAN5i/rfiYChAUl2k0yWfMhDEyax8KlhibDxmjV7ec/YI0FIAhoyKPD6kpnV
g3bXQm73UsjI/yJYoQm3zez1Sz6iWTH9O1BvRDMfvGEg2NMd7OPKQqxDWFPeM+6Na7a8Rj88/0zh
LjO5618KBTSnwqMjoVR8iXUe/ltfMm5GzQCE4LsdBUw/0nv4ZFwsv8tSadvDuLwSkUgJFiXVzSFE
b1g2uiuOOLrPS0GrfhZn140Bwoqk3fb7SszvckNnK1nZ9ULnKvxwna3WngwF+46U2JMHSjkz5b6R
fAJDK4EfZA0Sv1qa43NnFPP9Wcw+R1M8Gxwa+FAva/BU2IFhxFdgOwU9zZf7mvpfyiiCBDaYcnwn
yfA99/hXg4LIZ1GHH7OWUZzsIOxeY9+YpzFf0pUP45ptr/XTrHCqEuY+7CltQ2iOAHAmK3VRuT7h
heRIwPUpWDIwMI28dcJkhPcWrZ/525yYisP3gxoCEvWRGGHW0WO408WFQSeet56auu1Nc2K/4Wpi
JmC/ei8ahopL6Mc7NK3o9mPdjiwchTLg/ZJoqzgrwcn5j05hlB9Gto9Y03JA/fdS7rBZ04UWeFVf
Ntw3i1BUReT6DbM87Q3fVVXBjqEoaiPAM1CNlBgp+ofuROi2Pg7PtzsNA3qcz9z9WaBNRlKmGFiN
GVK7qlod97tABt792Y1szt+kUgJsuJZLMXe4RC7GADOqrOItKy63XtMRf4SkQNiIc5/gklha4vYh
p9DBfhK7JJV+OwiWJFTAq0KVwM2VeGpnIiPKuwaxdzmv88Zw9TpCnBEey3G3vyKZMlOReR28HXq9
gzY1BBqgfx/FknscElEimUm2qT4bNZYjuoCXtAkkrYJzzMyTyJWcrkq/u1APZEVZVPEqSPei6HiD
n9U0m7p3pOVUL3YJyf882Gx5ABI8js0ZTVl0Tf7JTMg7LQV3GfghyN/2SIQlVlzXE0muK4HVyX3S
N6kxsnBpfYZl85NOfVTBGlZXAyob8EouLtpcMZOQpwPXECVUt9TKaha0/kBb7hfwdzlgoZKsWtln
P73p3YTAriYerEGi3VhCm5hQlHzzhhSWYN05OummfjzIw6180zmpF9LXHAeivYbaltCTFhDitN8p
t7yAFU5p58ZrnxM3YD/92yNBvHpxOxv24EeJ3rtM87lJY77fJwzA6DMmaAjTwgHw+FGiSpHgiLaP
GRFnyhWLUJX1ukeAOb7ikxTjgslZHwTzS3du60hgRVmjUcVq5sePnnSucs7aetl5LbaW3bGDgrZz
u7CnASalgl1/6HT5eZpucHIOC7MfWNpDBzFcVDV0GXB3NSXhNgCSqWt/Kj6TqMsthZdxqRZlz+I8
wG9anhKOhZnInpWEvNB/fPMjli/vp+N2THlUoSr2s+a8cjuxulQPLanvEnQ0sDUlis/YJKoMrMmD
cTIgD1BA7upLYC5FZrqf368zti2u1TP3G0mAUzLjKUmukHHmUNmyNJ9f9TvkmK8ybqH8+H9PohSZ
odxDspEnqlMBtBDDdsSZpAs2afnneaayjiS3QkM6X2qJAVcZdyJRM6oa6+L3E1973A9VRSUbygv7
yzbyrE64V4A7nH3E8EapVv4QYpT3OEPheKd3HbFm7sBW68A9aHhVHl8pUXyHCmms3GGLUUS2Sgrm
9xfMSyRkfrG59M+hAMO1TJzQx164QDpsHiWkhepMPOnZj7lL2YVod22jPKptSzV8pPHqfdl3xQcc
xiX+xcw+fzEMnpGUe0a0LCJbWUPDnXmAJS8KwhAPtt3Td0mLLdslhFD6nWVjDsTxsGxCN/qYtSvv
53kQSjJPpJcajukvYdG+opMqB7YyFo0RmzNE+8QDSeCx2ZmdBqpb8ulY/4E9DlIDiXIncHU8h3D4
eL6xg4isY33Vojy+iL3KyMdEqvwM4fCM3Z5sM3Ghgx2C68WvIitlTFJl4lfTVb0JJUCZgmLVXjq6
3Z3lui9q6FZPneuSgtkF7EbZCCXPnnmW/VgHh9tkT+DWETNpniy3UBq5IKuwZCDtTkgLJW9zg1Ln
Zo5eEdtlx0bT/3iJK5KT1jQhd4ZUA5ppFFtOmBGzl37ATjhbF02pxvnY3jUQpthUJpbldW0/QjNO
OP5uKvenka3FseCZWpEVtKXldkEwtzZXXG2jiMHn9xm43jz3HRyLjJTnzdosGqzFLoPJlmRBQKpX
pzTJ4H56noouIw5mJoe+8L4h+oYJUoOMZpI/zpLh57teZspnIDQnEX+FR35p3IWqWLwmBkjgpRWY
tegqccNDyiI41jLmUDNIvL6CWVisVcirXwSlBcpIwEQ67is3txcZHxjwhjlzW+i9bKev50UGQ83Q
so1NpbCCWjYxweVJVv70OTZWJNoEelYcNWgPMyqI/zzGye8p2SS4PxvxwLy6x6yhrUSzKp8aE3pg
/UmAMoxjLp+SoAAvmFSwWGHnHu4/lEgpLBk4o51jIQlShWOSN2zo0wL6JEdEbJwtvgmzDgQZyJmp
VvyZYqhlgL8367aa4G5NCG9Zu3uHtP25XAbAWg4o0aUWuaWo3dXsbWC12y/SO7QAN4E8KtRnD9XT
AupOWKi2RVcPhLyAO0dEn50d6xqaHMTv99KFJmXEpg15mQq+zl34hbKrtjRKnboRTDL7yI5eImSv
SjDZDAJud1rilT/ut+w+NBpGhagiIjJ5tc2v2RAnMlPeDWc2Io1l3ljykMbBVI+y4t0N+EGjgwbB
xC1kxRM7WSUxb2x/blPkHbzHwJNiWg3dSCPhbqx9fCtYqU+A9J7f1HUOU70/COHD8sd391lZgGrb
bADaaOrrrCfmrxCIklk3AJJjsfNPTd5+apNsv+1rYa4iD0UH2KwEpp9bknr7meo6Gr1VrtvSqz90
NR4q6fyFdW1NMQGV7csoooe856gY3V83tQEC7/mn1zsJt/qv+63NfqrRQY0s2274FkEcSJ3jjjrc
MEIeBQhvNAM1IsuZdx51X5CrnGTsjfBvamj2IJhldGAwC1YY6a4NW3ZQULLqf4K/7iJQ6eZDbtkV
+SAmU+7KvRo7uTrOfJm0LzfYeCeT+RCdnHYJ1wej8FQ+qfrDVlx5DXiQ5GxJZ75+GahCg8wXNXZ1
TE5xBtGg/c+7MmvUGus3HO56WKgcoa4ok02GhLYjmNlzpbNrLoxWK3rbbnqibBMq1Oqv83ox7o/U
n7oxBi2W7CAiIYxh1yg/raGpaxr0/Y2Ubh3RymDBRLyi9Asqjk3foNLLEIGHEFef03NEh8ksHPka
/4tsRqO2UOcKOD7S3w8lIPYX8IHoV61Rrn5EJSjAqmXxbI1T8CNzx/AvlzQYVHVxE3yTSH7PYGW6
5oGbn8+UZPDUxYla5wNbZxuUwgNS9jtjPb2MEej/OHAk30bTQ80uZX5LmkUjjx/o82t/W5DC5yUT
2Byzt/P4M5JWrKJ31edPmNX7ZADA0S6N9JcyfpAFrp1oYeTa8+T5venbdW9XtBq7i52mUL2/KTfg
JWfn3MtGpCNt4Sw2BzohQv4vi7mnIretgIH+JAtqPJ+CGBbEJ6F9RBfITFmv1IvEADaBO81I36F0
//5OuKeAMCtfrLYL6VrSXA7oFfV14+hbhO+OBihvdNZm/Q5VMAvDplJvZ3SCaEitx6pyflAp/nIL
QwFpT0MUtGCGvrlJQk6ORNVbbn9kNIYPmLrqj6WkblHniu2hdANDDLVTVzKRRR+C5V7WVJmJW01b
Z2PIkaelmJl7rD7Tb/rC6LEswZTZjc84HqUZhHhLslpm1KzFfjrhjRhKG9kQr49vX9U+7r/T97Rv
RkDzVe/NK+sM5ybJf/hp46Qo2rJ1esnFXMya+TEpkLu04BlRP/7UqnEkpM76692areNuctrj2+sz
MLHvLEMEOfuTBbuNQlkTQFcWHn0c8jWfFIF4tFx1zAcm86mKoDmI9TIs58zuTrsw8k6sqOH3BlOA
oAg29hZQnP+Hg+1p/1zbAejCaEL9ohwPWjE1Frnu1nowVDjcdcWc5/ak/ejM6WLQLtAWPfoBDTFc
okZWpxxBRH2pgpOIbDjQL7ES4uUsyi8Gn2G8Wtaerps5nu1Z63Ft7GS6Y5oC7tvfz6sH2irZbtli
y5pjM5qC4vbW8JeGVpXW0Vb39ktfEQ1iZ6jDr89r8TrFGcT5mV46u4hpn94BUPK8EwFIQo9AwvCJ
tSC6mWsR2AzgpHS2f0UeoaEtuRqYrrBKA6cSF45R2nmlH/GINVw+U9hzXvvwov8jthgoYRzogw0m
MsYoSi8OF1JmXjXlhRQQQpC/O4NWZo+m84fPIC7p4nIW/BNcsQkQOfT4q741CswyJQ84P55v2EV5
s7e4q0O7Q6C11kfRNEPkAVecyBq4yoqkWZKUpXT548ydPJfUkjVotwKGpOjIXo8OVicKeQraBaIP
5LE6l5PGdVhbpaGLHegoVAZj3sQthwusB+Gc9X4sTSvB3M/6rHDDNJwXC9gepgAajCrX0h0tPu5F
EQQLWw5JsdIlijDd0b7rJzMawzbKuIFHT4e8yBGgLGqQpT9hRHdqKoIlZ80k0FZAN7IH7ZDAbcEs
K8cRErsDrWThuW+4ZcQGfeKMXBkJhcm81AfinCuf5owebBlc0VWy1x0dFp+ifejcZJmzM8JzfYbI
Xfi8ZmEpFZHgxC7ISlBUxmnUGJ6TdfHsYm3fjMpTW3yBUvqEihkNm2zMHY+sbYh8rgejVW03dGf6
JnI4FA7v3+hnowXUFHrDuHrKCil51E+IwJtROceKqJ7KQZNzDbU3/paYVzL6FyDBL0RSkC1bo/Ub
Ia+7ZzceKDloAAqi31Ic1pkuGwv+rKrNlFcEZCQerdSKGEoQCAKHPU8fawOwnvZGK2JfaxPxA3Ey
uutw79lAghwMFNoHi9e2LC+X/t/FUvrM4SrYBRZU4GCfaFav6crnf/uFQOYRZc/a0eF8tz9f2t/C
Cu6pZhiuTDl/pgtsOBJCArX3JRnxzV498hcEIAOA/ontJdVrtVStgAWFOKjUsxKF9EVfYROJ/oGm
4qryf0DYWaGZzJBLcgdvaAhIHBv5ZpGj+D+ayPHGMH+FGFxuWkn0j0WGlbKvBBPvb7TicKMmfUr9
YHFnX3f3kcuurAwLruXNne3ZaWib56TAVzVUs6LaOQb0cluJKyCf/Cw4KfKQgQchf0RZR3tKhEhO
HRdG5dnO9+ZeaFhvUAcxO2VWStNNxtUTZ7NytDzzGuDSDjmpQ0tJA750efVpYhZnM80FM6hCwnfB
7RJRlPwN96PxtFQv5gomA5H0Ul6j15CjcfloC9dXWvG39qJHN3cPXG1EfV2t0NunJweRWpkAa8MG
k5wtnLtrmF+ppUgvDdelXxMBtqS6naRHj3tEvq5Q+haQirW4I8F1SXqfRcfdKW9CzmxfXC5/3r0L
bI4D21cwFj6wI3tjJohI9gA79eUkyTSKurmaIlobqYLrNCmiVZ7OEif0vw1gJdmQeHCQtCJR/y7i
YBthQaCI5b8kspju4uw+uvUwL8BbdWgxt6GE1dV4SDkdwqEvj/Rdf2sVTxhcRfVuyRBsDc7cYxqt
qfGVK5b8RBTFEWfHUJWcYrQFf/CCzUOmBibQT9rW5cxwNFj8qne5A8DJpsYlngtsu8FWqLtGPfBm
Q9gOieEjBxPDk534YiwzgarvP4y1i29sh1zp11NTYz0zZ2OtMQbhxUEVpbGbMJpV6pJyXQAXCVId
2qByRyDpLp0fFP+fbxlp0tC2tVV2iZbNxAI3eyKLumih2e4p0VSHH3H4FmSy1yJ1DCoZ5c6kVXlu
YGHvOkYdFHRJq0llqNuxW1/TNFQF2BTb/aKn3TFSHuI1wsyAEd4tlA7vtjkXfzuGDRLtvlBAuC5h
uuJtVf046shc95gEcTNXwt7a97RUDwOL0sQp7XabK6a2iRIorjH1sqRoHEPX2rHBWXS4Fx+e6any
K84GixB3yTBTThIAy9UGqnxD0NRAP8Yi2dg5dtT1nnk/zTw1ZGohEhQ58DRUHNTDrXkI1fhCpKJ6
KyiJn4NACR2hWxo/SDT5OKY7btGlM8/5GMX1dBobkOtdUCBo3WbQ0ggWGFhoG/6+iNbMtcd2lgal
rRu/zENZSlO6eyJA7zghKzn3ikQF7DOr+NU8uUGUzazaCLtnPo1HTbsk0T+d9oi2rruOO+iLIYE3
Bl+9u+81kiKo8VfVYBFCaRFoLOvt+3NhTT6jR9kr0Fvvaezyrx6MPBXoeGzgrS9llYoBgEAva06K
xg1iopdHgp1OxLu+9p4sX27iLcEOoFDAK4EwT1fwpIjkUZ15y6Lu4BOqFk/rCHu+wZ+HHTHN82lE
BLlZ3VKS3iAUBIVa3eCxEsDgABagm8oMlBvmPYRW/lEbrKTbNDb1Ljz1SlKC/EsI61nUGOYlxfvP
v4hnd8wsKfBwD0kLD+9cXX6Ex9hEJwvYavlc/uWp8Ok0AV1eTVkeGIs4xieJussZZfGPAh4Yzbu+
ZvyI0Ll8Rx4juCIdynX5hKkI9pRHCi0rewfI4B7chjJu1dmcf+eHf1U/XtwkpEhW1Z3q5bQoPXfN
s2nAbOASScXRjy7qHXBayeN1IWWjNy78b649JT1A0T0gHZXTIke5+uNOeRVN2fLefQhFR5He0m2o
wI2cLPYKkFNYiNk28GfE8UNe3mvnTC/gG4W+99v0SNyrayzMRXDJhtBnBnEk8XxwjCCgpLdATqDx
vrnkPqDE/KZ4vXecwuTI7aNbNNZXHaZsRxeZ5KBgFeWmGmyC7+2Tf99a7iGxsyeh314BHztSIQIW
2BZAu29SVZWVkaEC4N7VPKuQRZpli5UxzceX8b/0oV8nyd6884VqbBCmwygfcQGB+yxwe5YAtoJS
7TAiBJXFsHJGlNJojSmkxJSOBAocxe4nQL0WXGZ4qTnZOQ59pCEoUIgs+uBFjfVEjWxF0Jh13LrF
OgbbvU4Fz5fdDc4igmcWM2Coo3Ce3zrSpQKfTngdAUPbjVdwSUxQjJHrBS6VaSo32ObsCSFaBRJw
OeTPUPEpIGrA3MACloD3HLKixhqDY7wDIlkBWXtIEeNP/gxmYTPoUePSuL5V16i2F9tCx/Zf3QqD
NtIXknc0YMyHfsTqx9STTy4GA8H4ebTl8EN8h8xcx63MH4WMkNJE0hq5+4ehOkE1X5yeFc0SXhNX
dQoPAZRozG4Y1Y6NcZlFhoX3cp4GfjZOAc7UoDeGng9/+LUuvpnhWRIomkCvEbPuO6+zLZEFCsu9
v1mHU6ZRVoTee/gB67S8JlJq3Z5IaGlTeij/xxczjP3fC1G5d/b3GJwe7jGbYZIk4i/ju/z8Iv/I
GNlP+M0aOeh2ZcDnCGI3ORYjO/72o3fTs3hb1FsG0j0cIk5L46zlqpYOCRzZaZpPsEns99pwiM0m
5DsJdw+vHcivNP0tqiAHFSwXTZLgODvLObJi7KWSElAngWuwZkhn1/tpQSPSoltWuMDBDogoSIMV
M1wOaHgI+TBSDdLZlOekfpOwpi50zFVnCXayCHeDbyVDaIzhGv1GfUixymXTeOr2I/f+af8KPZtl
iGzIKE7iuHCbBcaB6ZKeWT1yKvAM9D1Bn58DhM0JjLShkkw21i1OQoJOJUcen+tzjQH94/tMlASw
4qUAUkXj3YdWrOPDY/VhZnm98wH7Rwpb24748vsv2EueqIh1D369dAZDxBYIBp8bbOSYh81mgILk
ieSSkQQuCeKoCMM+pog8FF80g72O//IFloTMXyeEPvSR+2lbdiaWOq2m+td3enh7nzuscOv/5h96
j1FxQT87+jGvVG7vxEQtf+XyYJ7EBGG4VdLuE4zhjpv1MKyrcaDYKSVTaaLN2gBrO3DptOLJs6TG
qQ3L+NUpqbHcG3xbl6TWvzyL7sHacjjtFCtPIV++hupwJvBV8dDn+/Vv6v1BUZgDFyFCPoTiLM6p
EsFLbCIczwZJcn6jfS+SjJNBmiF62hoI+Eoruat0HwODaCk5/+hPogtErqQsMKOpzIw0176Y7CnT
V+KqDtVBwcxd69xMmurfuFrdUaZLGBn30TR0jrxMjIV+5VpPNdyyPfwvVjDoonm9XMr6gSW+1lBK
tDsJhIiw1gNadEXXKoQ0T9yTePvn0UY8J5/qSbGiFCvnLNi9ZV/u5+qrELvsKE2YRpPxUDBPCOrV
Yjdo3VgSPaf4YzwZrxnxHnR/u/OloraL3qB465cPVCu2ctzAIU4JMnEJ6Zd1EvHNo0ENIZRQlzWp
o/Dq1UR3gp9ZwSanA9dJU/aFNeNCDIHTlDvxOs9Rr2szCELLBiy6HPBa6DBvUVlYTmzFH4Sru+Pw
wIK+klwNdsgKtNlEPy9esp9gYNWftea6za/58pqouhDhlMRae7C+O1AIpxVXHSghdB9yB2RALDsc
iH95dhkW8tukEH0PnoooG+M93bJFXeUz6JBAfXxzMUgoogn2EBmOEm3QlYQPkHBLjNVkhKhF9paw
rqwQU6qiQg8wrcdRmCA7nWRuYhlnYjOS8fMlJ1tiM2a3oQy4Gbzp33txixSIer58fbfMWxWK2IWW
O9QVUsIkdhKZb2RUmSo7YcjbhvcEcnCo+MXPir3ZG6RSc7nAy0K4O8FGJK0XPSUH0AcTYFLypZKM
E7gdzpPTWTXFJV2Yom3M9heXEh6fTwyP6htV+n+vKZU081h1+HDh++hxlYVk10jmffhSt1u9ARxu
AaCXTzylIvfM3IVzJHZx7RYadp04gSLoQTv948gz/SSp30XiCJJ+sSsx338jrd+4m/z5JDhxTTID
atZlnVV5D+ePgt3Ew3LNbJ+JVxWcV889i0MX4q5Gry/U+vgvobxQSUBHWTCQcRZ0GJ3Dws2lUWvl
p0WKXU3RhGELySyf+ka2tV/pWcJKztB1M/Azy5Xj7MwRCHoLbcRg6k34uSf0gVlo7L41tCzk97I+
hhHSqS242IlOu6zLeX1lvWaMzA2LPYQ1SSXbdgtYTVMi0j/z0ORpwd2iRxgEKcDTRqh3AheC0KKo
LE1TW0J4b/O4ShY4wcPTFH5WN1nI6eY2Zjl3fZW+ZIaItqFrQoBrrvwLg+XCcVWr/FCuj2lG1eFs
sS/t87IDCB8SvVrdeNTsGmKJSqKxUOLLW+7XoQ+lBuHE595VpwvV0eYq8QFJwxQHnX/3eRCxqJF2
k37RmVmM44msM4A2OhXfNGieNsobGIIbc6ZGMHwCUTwKerqjtY/0HeCLjotTS9DY3Ixgmz7akZx3
GVrMfGYM6eMD5A10RTJAnw1a4gK3Mccc97JZdmMaf3g7HmmH0RaQ4yhTzRH9MLGc/UuZcYocp2EZ
kzn8ZxnaafqB29u2agFmIkRxgZ5vGzwU/ODFl9Pj6zH0qkxg8cmyqxx4+5o7yA1bDf8lS29egsvX
vQ3sxi82ehbMWT4cit4Z8qyecT5jnATP/uwCk+JlwYgXB3RGczPsd4VKUJczKXRDhAf7FMlm0lE2
+0NTyn4enhh2Ig2Nj1eP794KyHhdGlbl6Z72rO11fdVRoNc6OL71iYsKnSnCx9J7DWVuSAEHiPbe
HX4UjVF1aDpuKBfpm1Up5FreA7XI6u82px5pjT9yJniKWNaTP1m+OWpP9l3RTdXVAuJx/3zis5yl
abQNOB6vcQv6dEeHdtFVaSLK+MSx9VD1mxXUspOROA8Y0z3rz9bHaaxlfG+TU2a9uNCiwMW+Bkho
MNC9Q8Xxhh/G+qSmRh25MEedH5SB0O1ChkzWFxuG1Ke0t+sXaAlcwwfpCMMvR6A5BBd8zQ7nrUOH
yXaMefH+OuPKEhYpdv+b85y9IDxTNB4aQ9XaLegx9ZAxVmWYOuL9US47B5NnhdT88lAm3g+NOdBT
WSUeUVLzCXkZ2NcCdTy8Mc8gPoJMkBj3P4MqDXSx5hir80jiKKVwV12k1GJg6XUNPbmL+vL131lB
vOhD8h7aMU42XUavxN7EkgY8M2gnPdPX4hx63kBrOvPveO+2Hiu1G2OMBRWPhtDMU4sTiiGMgBUo
ZVx3GuKTWptRWxSUe4/QSHaBhbgxpQ9cT8vDhpx4/Gbd5CKfOOmsIjmXb8bnimkkq5pT/Fxd7ptl
13aIsW8itAXWNbVCGhx5mYT0VvQMciTZkdFm3oODbYSIEbgcOZ5u5GHoHRoqZgEf9Rx/BlD45ZSR
wJ99YYNGsyOc9LyAPOqqyLeQn/z6Km4gEr8HCmyTAIyeEg+/kR7iyMHPJgtCs5c1ZTmdubK2a38V
EYSeIk6fv/Xv0nG66DRhtwHXKpIBFA2l/q+ZnoASz9l73n+nPlZIKijtFajOz44MpcDGskJFHdEr
pYmH/yeoerwZg7GXo/wsPulOP9UPbd59zrCbzJKj5d8MbUeVKbIBjhL1Kpb1/XRR92yAMiIOSKX4
9ypTfBt5M8zgRH2jgwoaAhFJYrvTxXKZFlcZYAz0ZOX1N6OGQ9kdO1wPYEyxHdEKndB+Rz+lwprB
yT30vNhegaMeilDBXQcGHGdtseIjPI5MkToIrfFv8ESJscHzvQC65V8R9j38JSmkhXl9PaNi7WPo
hoXjJlo+O838TuYMf6dqVQazzy6f0rXfuIe3xD8Flbvbfvg9wUlon+L9lQsNLdAUQQWx9wNrwH3e
y8+uDDZo6n9vQInM+h0uFJb+FBDykFvbrnlK800C8+KeZLoyOf3mESpozM2qRXH0WdcaTpWnhfrV
5f924PiwriRBO03bJmmNRIoMBIDYSLUmMorJRfJCQgFWf7R/2koxfMeYfve+A3xQ/96UEjF12UaS
NrZivGCdY7D4BEO+oX+p8KKUDukldkAXqyu3NrKUBXVCmGWXhm5OZd2UT6McDd5eUxAMHHcwaFuI
SDQISWYEOuBbHlfPhCsL6OIuZ3eI7pgKPcVZLbxWZokKhsM1G8zao7kMtYHD5tRM/XyMC6IlU1sA
qiL6InutHfDEFaIlBujyIL2RKqLUhZJMgDKHjOfQrxB261sU9j4QfCNzyJU8HtrYJli6Pqz/6Cuq
EMib6I0x1Mc3u3sJyKF9erKxF4C9IP53NSWfcRcbB8veCRbp8t793Ju3N00R3fZ96iLQ+c3IZN6Y
gvMNBxo1ypLj3dexI/+bnx4XBgE1HVsnILg+phIztLr8Pzc+ABc5mNLSqlBZ7gG9Rgr/mJoqQVeP
wkKmWKKEHb4fMHWmkP9Ax5/7Cj8UpGCwF2rpsKCsrIQf71RsBhE8d2LRaD5Pj0Yi2GtA4ue90iU9
eGBfx6AQX/tUiVtTDR33eYLe7L26DSQnpeNMjde9MDAcLFslrea7QYFIa20hlpsN2nAq6lT2Lgo7
B+tGcVnjH0vgLDyg/UDsFXin+PDGQvey5jE4Bv0806Mpo/nTTvJnaLLBD2seMNHWM/rWpdzXXZMl
w42VXXHyZEgXuHCs0an3IEJvhzITSJS/Ix/8S/IR6jSk97sX8aE1c/p6F5RwkWqckyMARydw9vBb
s4uWuvPdgZH6VIQtIv5NI+linzBIeHL9tcsoNtKFu2C5L3j2sqzE6t2KIV0VQVYMRxB5HglZi/50
E2Q9UyF1lHfxJV5C3J7324wa2RMKrTELL44X6O5zkgXzFi9OBg6lROxw+GcPUM+OB4M3H+lSYRbD
Y2CcenVwsATlypsnue02MxMZt/MBTPYTJuNmYbRYpIgwV+YZ3QdxVFh8jbQH7qcmWlwgt4hRKl52
iZFXldDbfEvap6+Gt893ofoCY/7NoDdk2FBqZ3YBnHyRuYl+/yAQ49WZRRPaPX2GGmOG3AZiX/3J
Mf1uxgXBAMFM9BQjTKycwC0eBbXgUZ/3ocGzYA5IQDY0mNCdplL/R1Ujbc3rIrCoJbCzgBlrQXBV
IjhOEgAgZQJeVR9QpnLrN1cOcmc7sEUIBslPGZh3FDuPUV3tR2NsTqV0XbI7LZNybx42ZhFgAgQK
bGY3rcFxKFu/qR8+yNv4e1NoWULNCED/eugHBwvpuCtAAWRIDZwuI5Cfk1kxfBvZoNtsOLmbF+Ey
kMw7SZN8L2/5KqK5Zo2v/r6KPrtrFde79plehEg3Y2qIKLipWJGzMRATtzccS3l8Tw8/tKZy5MNm
ty9wuLFE4IUdJGKj8brvVNKK903+NmEGV54RIXtL8JVuJZ0RXgFgjMtNirVSJUCqXFrq1JajX+vH
6AMa964e6KFJhHsbYHEBWDWdzmLRjpOZrAkj8yGkg5VOivsNco2ak7ERszWuBhoEYJP2RD9ENGj6
ZL4c98J85IvLXQdVsa0buC+T9iVsY1mRq4S4wEWfzLW0HzhUumRaBybsMex9NJj+MPnxAHqZ8PFd
LtidoHtTMz4zpgAEJJ2VSD7MEwdoY/fuM2TOOxz//sqvii5fAXzVHyXOXJHe8nO2+iTDIwPo3Dv3
HBiha1pcmb0xaD+AfN32/DXMxOlSR0mcB+wQdfAejCJVzX9y6HOzlEQm4GacVpnBMzPwfV9gnWnH
pm96VN4PQms+jznitnTpP08HoYrCu2hzKmOLSy/xzCOKqPLY42ct9VnfW5eBRLovOa8WsB9fCMrx
X7BHDH0jK232TOPcYBCy0eUx9KnWHZ83oJAFVfXH7m+gmwiGfHDo1Pn634tF2G+6S0RbPG3ER3Ke
tZ+4+oW0egeW00Cm59OJS8Y2GQS/1UzHiNUULqLDxqgJxA4s7kTBqNYuY8UjQ5SNglpDBWtS7gTl
Z3y4f/BllpI6bINIy6pnCNphgGjeYqC+KV++D9O6M50zwoyBQFiE88XXZFJZJ4qyJcvlSiuhrkE7
N/lvAEfUbtQ+fw3Gn1CU3QweyVng8dL1Cz7sW8ilr7tgyG3QqdsAntV6Jbot0cfucN7VE9hnjyvN
10pNmd6ZuD0+32S1Xqi+T2d/a4ru831ZIED4F+zfkFivouBEK+wecMNDXmPrIeCSuPz0Zx3MClAa
/DaZMQIglcP3nejngcvDxGDCMZHK+VyRQVSA6lpiLFR4UHMkVNbnDwSluHfWR6QpAXa+9EdrsEfC
qCHvNQ5zgP9ploWj5G9RXaFU7hjhBdIxvdJvb92i2iNo/Z88oyfhw7KT0PNn+UshtM5EwpUcKyx1
JwmnlLb7gMa1PsTzni0S5/Tt/+Q4NBYcDW54EKB2OWq9LxSyJYsAFOz96enYBdS/V48ibXPQn9AT
ANxGaFljwEaRnL6D8by3DplhhRRTDG0wzVAUYG8MpxVdaj/O89RFwHVy3eF/W2Kq9ucPagw+W+Xp
jYWPeryfYImGQS+udTTiohIc7BADaTKlyVXF3SVW5oVK5qIejPrUJ3p0xXitCjOacT4djtrUkzRy
OgMH/I6KEGExZMm87hZoIj2OkYwAc+x3P2a2yIv4IUR2rtkuXbUoEUs2AlnHjla/jiyv/kMI1vJC
3NYTzO7ThMsCteD1mjDre+wqjI7RN5qDs6N04Z3ATuXlN43Hkha2MBvOFm2NXr9iaYui3waQyXoE
yaLxFmMPSGDLR5ajf1BPzrSnXknX9TqFHG4Vo1O/q3Mnxi7wyGRjvnQAR7Jlvvm8NX6q1e+nZRe6
dDPr2R8n7UiVtko94rt/d5/h90VVl9Hq2LSAvLfVFWqj55DoEof7XnwbK519ZV5/SuGtAFZBhLeN
5EViT7sv1BlRE03HnzQruYxH6mdni+ylytEFdySoE+UQF8VK3lDLBq3YCJR7/lt94Nk0EsjAepBY
RcScf07sHvCOYL5MeLTpJZmqH8XJjktJh+unvzcOYmA0J7TaYgYAfMwZJJ4WRJxeQb8hoJjDEbDO
c9h5vBchSAOSOH9/FH1ikVzcc+iGfrNtevc48pB2Q+xYEsBrtt5kVr9nk5KUBOTpPqiEkpLC+wR6
jp/RxVQEKg+Fk4a1Jtp32CG80tyVPSyz5KQFW45hgjIoej6a10ZNa0cRK2QXoCO47XyVuksE3UZe
0hUl0q253tsgKFG52oK20DDimrRKnq1AWMvjlXu/dZwl/1bXsTwt1AqMPqmImLbs2MxjUE9nb/6U
lemqlGNsRZ6eo/PG9yNWLxq600vAaUvE5y+gviPmTfOKvtQaC+juyT0Xf/P6oJt17FgZ90CJNzDu
q7Dy2dB/8OEHH9XSy1/cFfGensEaeBxCH6Zcsy8IdjtG+ok8M+T4ByPjqak29Oapr8P52isVhLgJ
9aVnscr2NKtFI8oPBD8Qb//wgwGIELAxaMIiPeEN/N13FdUpiJ+9ZHNJCwYdL1maAd+Z/nhGVMsd
TkQyaq6nPJFWClH9IVn9Tw0QqMjuQb3b1O0bcAfUiSynx4zp49/Pg+teRJ3S0FMDDeol3JVgcY3K
v+I93V9pSOVvzh+jpNRPElaDbJif68OCINdeXZXgANpUijsgWaqRbZv4/yesQ/hCl1mStN3gF7fG
qa6cR9tt15Do61onyFK5EJ7Dh/piWrUNYH4qOAqAeVRVsHbR2EYkA/UeBlU3YXmdZ26RZXgBZVAe
wIYvvPVG+NNbAhe1AtDn0hA6+cgyvVGugYkYJgBVZQoKnGBj14egcIhVV7qkC+PugGmu8NpU9F/R
jt3LlzLHxRr3GYDg55IiztHkMXUfAOBdzei7MJCDtsG+iVRd8EyKCsRbSsAAnMm7M+iJsMWpvCwM
YbmvPo2+9NzmdxE9wIJdm3SOZhJt/ClPA5ilR/MHeXx+YVGg55+qUP94oDkIgbIkIMcN1SxUkhmc
xoylPluk+yQXHiQoSpE1WEZUO7O8g22Tnpb1utnWh9ZMrFtWLUYlNjhx3crjcCRHG+wHxrIxw1Jl
Vt0iHkIfUH10qLhDSe1JRnj6KgCBTDZrQWd5NV5Jy5FsJyDugOyuDO/rdmGc57I9GHKyJhS10L0t
ozPfs5sJY2GsjavzrVNB3KDixSlGN19Nz6Ao8n6QfgAXOx+e8ZRWXNObBbSgm0t4QXqOsFldlMIU
XiFU701N2ifpVn4o6mqq+YbaCiuNKESCOhJ9+AZXE8pKP215UeVfHvuNiedXUmsoVX4PnpezHBrz
PNldYfi4K4IZFATkWdxlXdY8uNjnHPl4REVkQPIyTVUO3zRzzgrUqGs8YNcuAsCdQ0pmlRNqxpQO
3LSB0hr0PcS2LmQeig9kkdnj8VxEmjV8uP33V8bmadFQsUcWNlvbNvUrHmUffergQs5bLfu2e637
CxEbmNt3qFiSdFSyzKOFcvCdXXYWxAAbjNl+1zqTCejwjYpprmnGvJ7cAIOosRiMVDWrHEpUZ5bn
5dHVOQFhqIKPnESF+Lm7kpxKL9iOxXk2OAx9GUoJw38URyDQSLB+6KWaMCeQIU7BqGME4iXjaVEC
9RfoEOfyCH3mRJi5Jlw6UC/7LaC8R7s7XTSM5In3ZCJIxXjBW3Dcej//HxSJ8cj5eJskE89abnTS
+zyNcqu0K+pAf2QZ80s6G5ZYWxft9izfW7prGqRXzSvcP64BksbbJMWRmSkbM24wa6iEUDdV/wGB
SdES+bg5AW4CFxRLyIFxVV43xGc4zQFqm8CpQIYx65NOT7nNFMv/0ywOdMtcKsiZ0ZHtNzq7WnV0
sZhNE5yNylwIjVYgNFt2/WTlWGVm3tzyeR+KzTErke3r8CgEAy3aAmhLELvnUYULEHatBFbnUSUP
mSLbLQi4QW1hWQYKprRMQZxXMD23uQrsAgbURHWSbBwm0arh2qWC5JIrsI767gtmofMQecwF0paO
uTfbhDh6tpX+FQdXXtCxlzpEK+BVI3DGbp8LLre8FTccYVQMJ0B/41/QSfP/389Fl69iHrNyQnci
jXiFxwQAHc0a202GCQacbwf2gxTVw9aB/tkCzADTj7dacBVCZNfHnKCm/SPV5aYrBAPmKB8VSbIl
GR9UbWhpNnQCAKrm3W5ghrWVVQb1FNeURXy5p7qhDd2ZrI6wSRib1fRXrs4W1RfNmduGws8I+p4J
L/AqsWAG0FmV6TUaIBYbCm8Ynl+4GrlTnSLgod/7HbG4vBywiZfOhI+B938cSFs5PLsd1pmG9DvH
EykA4tIMgUmzy/K0y3T5ZnB0+p2CiOqBZAtwwQ90yiJG8rgegdbS5PAfD2PXWZ4wmCpY9Orp9W4/
SXAzz4ElTmhhd1qnTo9KZr5LYirUfKb13E9N2Kxoi6qvIEs+WKcpiBTLmXeK+14M28U7kUnZTt9K
f49q4BRCuURBCGFSovJtBczixudefrGnr44OuW71rTLgIYteSgUMF46haSInZtxvnUVQbsQzOpEo
atb1LC9AThuvnQ3VGHATnBDPu5cYuIiVBPKi66NHS7zCNhGs4GufeorVLrx4zBy5LRb6VFHbt1I3
/1YV8ofCOV+OlLMFgMZlpuasr7LtGYh/+OBrL9ElBcy2/hYdXlyLGVDaBJuVEVEYM5JVTYSLnmzf
4PS/fZgghJcVbTREf3DT8SZcWkm1MFTcghG+gVZ//uOau1pJeimnDNZM8Isw0m/uSDBrbvEztDMh
Q0UA/7ITH2QcFTae5SVXry+Jz/CfiZbXHQ3JOag7l6WuSbhoPtXyNcy+qr3WQfNiKXOzUS7JyUL/
PUbgBjm7wYgCj5TJ75gGe7t+5p1Z8Pe45bFzanj+rumhsRFwIhpzdiaEAE5W1Tgz8OyzkJJARa2a
Hyjtzd5nSRpKUcwwJyv6ThzDVikm7W1kpckC/XOzX08wVZ6pWyBkmv7DnlOi3KUEDairb3rRLQpa
JjM75u9YREErmf1Ig61r2KRa3eVCly+OsezGTqGRC+fAyPsyY99SFDQg+qfrUpg646rhpKoXsfv+
A/6KF0YtliWbPPrJxQ1szc6+Ozcv/j+wac9EwxtAndV7Uwo1ItqcuNlhhMsi+mifnVbt7rYygiIV
xjMqLiCKN5ZbTNU6JCv39YdbP9e7mp/e5o/TuUIwxrDXeYVPHTiCwV77/Yazb+rKL3Rw6MIP0qqA
uEvry8hR2I8Msq53+38mFZFnfQtxSbvkEbPikbJLlMzyCHN+0fwd66558kVss9cEtjWg+fx03gui
84xmmhi63uZ2jmFTRl4EFVwArgeXMBenpMwfB/PAoCmEKiSBYEPvsgGVSfsf/Spjj0BR9XwIgzsu
H0fLuGjpeqJEA1Y3t45AEH+uN9d2wClz0zJXyWGEK6GZug+uF8CDl5uyGYcGVxNiUlSHZRwTo7m8
tSOtFavK2Ii94STb/8kH45/pmXPW0cfZPfOzDqsSDMRTjErLriuA0Iza+/Fdxd/my87W6YAnSKdJ
TgFYZAGOebtqrEZqgCqYotz4ZDFm5aT0SNNa01t0X80cuTydxOLnOVn2HjzDjxwIs8OElDVykUIy
rD+vLAOciCJkMmcYDq00wW1NkSuAnAQLhXq9AKUqliNW/GKZZjzHwTyhlvsphwzvhij8OKHhUWQX
OAGcXUzC8zRjJoOGqiD7AXi2GzU0sayZpuDb2bbzZyVw7qoEx18j9dPhn2Ncd4cGA0ye/VEppsKW
oWlBR0ge/9dtSR0bMR/wnyh5SGvpi+IKDpYmfc7dUFu7gJWgymYkaSu8hzpaVWafC6GmGJ8H4PwU
iR1CJ1QxTU2slrvfUvQdgh8Rewj5lSl+9yqQrer453nWcnOGbUt4Z3gMRSuTxjjXsrxMK9GoFMZV
uWNTEwfzYlE+nt6TEV74+MXxYBxtVJEhV8Y6iaUM/QdEo3Sc2q3kBVRucx9xp+gGgSJQNauGp1DF
wLi69ESpRhJMycyq95kD0+BREh4FfZ1+ZdS5Ip/nRXosaVD5VNa0VpqPGyQs0dJyQPNVgnEi1GHo
tS4bP8gSPPsOCLPjsW3cgrA7QOc2y2hRaQy9dxxMl6diaLip2A0ElsLdlt44wQvouuGv9/YtY9Ne
Sr0zJ2ToXN5BkAL0a2wKovHyyl1rbnlWRW1PYx31Bg6v+ge7kFmOz9YWd919y8X2G1I8bWB3Q+BQ
8HkRbh5Ud+GmfUmBKoi96YXgzAvWa/zzf1dGj2PEHgiDXzqvI9TK0/Tlg4YVrApYo9RKhtHBmtYS
ZIQtQinCunVZgqHGZIm6UfqzaVyEplQRh9rcsvtz2kp/Df4NY2QVMwQljvHiAoTNzrKd33yze4GI
5X51wGkf63KwizHe/K7G/VJSIQKDDjebWhe1VQpenTwKXvqbvTHVFU9sIgotVRA1NjVVJRsflBaf
0ErFffUlSRj3BFvI8RRtipfsMD/rQuCrpcnD+fq+macbOjWmy6M3SbG6P7zUsWVy3OwP7nzD1Gz1
0TfoEqjWgevrpkDnHw1E6Bxyl/21ieIyVUxeH3WYbHLz+SfzhJREohN6HT9ZbhvYPtJ7IPqPbY1l
4wJqSMsoKl8ukZvlbhGhRv4lANmghcg9ehSTrxLihpje7NFY8xbUMutT+c8VLyNTWE420jF206AD
6/pCkbAiq75Vj0hTr5Zb9kzz+Qid7kDF9VS/etvwmh1NiFHqQS0bUfcWt5pbRh4Tk1BtD/B5WFI+
+whePky3WUvepSBXaZMlkUw0LVp2uFB4U6KCsTqsXx7iRVdqixEVqzmltR6h4Btegbs7t2oo5K9R
8HmflhvSyF7qHfBM8LlR6JqMsoFd9c5fefibPebDkY1SMwo/qQ7nL0p2ORbPoZX/rrH4I0cUqzLN
U9+GVoeiDldp5FjgpwaSRJ2pmfX9bc8DIzQAxDo9ggbKzCKmo+7l04vOuGsxpiU7yKXg91XbKv9b
m0pmsuWKTyl7PmPtfsCWgMPDuTzKGee1DYsNUWQpUY68fFoHTBnAD/KJmjWBYM3ije0znAHV3BlZ
BgDPZGItpQnaEryUV87Ab+foa0UvudTKVaUeQnsYL1fOGBm8nqlkM4aZX/uCAg9hlRSkI57EKCuO
4eyUqoYeiau46+FMXtQmAVHuye1ZD1O31ALbakHsvpU+hjCTealtkN4L9h+L36q0jMaRLjCEfj9i
AEFJ7Rko55L0CPOG/9dwWnvVvs0X8CGTqEa9Wqu1b8qSmfPjAUsmgaB3alC/ZLWxEAbS/YG/V4tx
PxgwMktnIl/Ys61L3X3sc1fNDRXBHcS28rstTUxVZxm+sNd1ERNU2fwfAV7mO4jhgildaEVMBI2d
M5oSz1+IncwqWrkJhw4DcDcx8u+adupLaV81K6Ecaquyt2c9FU9kd5AqvBHuucy4Q/hfxHP/X1hR
4PGxWVlPLsukBQAniGXr8Umw6o4LC44Kxk8JbE9msCWBxdFj4sN5XbYUMod45Og+H0uWY+odfOnk
UQ0dc3ISlwPLkf6nPvG474IWV/4p8QRboSmD1BMsDuMrHDYLkFjMOrypocRY5l/OkytgPfWGZEbc
vfkmN9+Ke5A3FfeA3BSouaLhYwECx8GzCCs7n72AAm1OwgxKdkwTa4bsOOqVR9FSOOKF2Tq704g4
CRe8/I0r53fHW32jAFY3bmdQt1cm8MO+HBGRblL+D54iAtJj5myyIG/JLlev/uc/Zn1CSq927VvI
Z1Cb2caHeFLHpAtOs6Kksr82K4WcOiKxmrj+ynjCwn0Dv6Itz910E+NYJ/bAZg//n0yhBpD2saSs
itzzAu8fVB1GojseHdzz1ERg4nzrF6D4oW4ZjVUWQyKbO6/ojjmqNaU2vVwM6QBOyEtvR4UbAp+B
zZoFkP6iywskUBUi4zYWBZCS3UXfkcLchfoo2NQE3XAUZSgWlLRDk8N5OGsq06HrybJ6wNDNdpLG
joWR9iDHp023NA+1iEwCds1PVkJ+SqEWuhjzYEB2yVcIT4L6AXFup4rV+V/6giQHr5TrJ2RyU65T
u4vlCHzk8nQAxH3xD3sxTlFhouo9Xqlui4MkLU4d13kU6Z4uuegZiPCFDV3pIFoKRlWIU7eFo6XT
AtWh35aGlQxwYyisKzTCo+/y4m8kezI2AhmlLzU14KpjXkVsEQenAwrQgvDwY4XIweX1zsQUCvwL
X8scttWEZjheCsheud6dxMMACOdkRFBqeOV1QIwA41T542gx5jxYcycGFttclY1R8TchNPbAUPZU
ahG6KumQ4PpgqblZb3R0OALpEV+fKa4EpOsqrrLNHVg8OZl410LkonhU/d2la0s5th/iDAhxw8Mb
+E67OJvEgTjcT6cefgRKB4TfeSVnqyOGNvXJ5Fjk8j7C3gB/ctwBbvjAJXA6dtgngmNzKevgYwio
x7YJVf3oHM7YYRI1jqjqKAHYiO1y6sCcbABTSPQ2UnEu63ZasH4t1xQvqSQja5/HpG1m9YVMRcDA
IIyyP3iNk5aOIFa7m/Bpdez+/Op4m9jM884E/GMCev6zfTnQjdqZuYJnh/DnXQp+ZRyTFAtYFOe2
vbQWRLEK9+QhD4AaQ2SurhXHHLRQUCZx1nVyOrJqGOIK3/gXEahUx2UafxR1O5/B2q7Ac/N+Te/Y
I28RS6o7p7+mT7DXS/5VM+cfSbjMZ0L1Zx/flSVhs5C8vDaJ1rwweJzx92Eh8wnYct3j/Zzdxg6F
n7J8yBPvvHpY4VQlbnJLB+iXdDjfC1ciHHhatYULmChv+h9+LVFs1TW80CiL/VXyOBp1mNncOreD
QJ2URYja8eHle+BAHx/l3VaSb1m/7GceOwusBLGu4GPPB98hr8AsiJGx7B1k2uJwNafisN0xyoMU
dm75Ajim4DbpPqVp2wtDl8FNspDd5tbptdakw2sB9SDM4w3Kt7xk/U+U5fItCGqvjVqqJyDA6ffl
LTNefivDbno7yrRK5tfXN6E8VLo8hG0x1ZM/cCmviObbLraEJ5RupbmWz7IBpP9Ak/XYFhyz5nc5
H6kFy/7EUtZS08MJlUQbykI/syvTHFgEqVj61VUqVKKs72+l8HjAeZZ6Ek2DgEmuJG7mf8+rGpSC
zvOE2KW2IOtisjuahSDb+lIvjuUleVyLG3+/82hOnc6jHoKMiwjhmS2SqtAz0hJJknZNcq/hm2mL
vObuQrP6mwvvXYdD4Lu5RlQ/d9P3aZm5tQjX6Xd+v0x+dOot5tWhDGSLIp7WBEVlid/AyzT9JCQ8
nK1GhhK6hO97QFYqE/OCYKaUBNGOeR6A16ACjjnEeROPLazaJB+yQIAWKLFu/2K6fS4E9QNtwvuK
axckRV+3BGdW8mlhI1vN3YQQl17tyxy6XClfKBnYEbTAQqVadXG5wuQ6RgcFfli0zEYZiv5/tKW1
HrA5MEL2ypHEuCOLfmCSwiWfNJpXS/AF4bdcNCdYdq7yB+hSADh/9UHfb35KyukNxn28wKTZ0QIn
DLfHRDgxHBv55S9kG7xCGgLMhN+7u5CcUARukXhRRfUzYYFi6TFiEI3SqWGqq3DTUGk+jQej3D4Q
aHrn/jqok4icn39BXiRY0xxnFa3lijCDGiHWDL0+DjL9SRr6KW96OLJ52HL3i5AF3JjezKHr9YyF
cjavBq+ybXn3p/qWPWOBRHTl6bCE01fsAmglmtqfWJnWHppJW6Ng90us832uhMzOWtHKCnZFULES
WvO1p6ojDBRLrVq1BIHYvk4Ra7jB4PFq4ZOHUnGfW2T1u8p9Xdlg4ffdjHvoMMvw9Ac/9DA+k+kG
wlR2BIuKsgG13TvGFDwFCh6anR0mrmphjbHF8hDErKX5m1TsJH2ZCl08apC6N+TAeR1iZP2FYaa1
3kJxz9WfVN9hvnyBUCFK70o5UjGe/9XNrq2zRUshqlXoJM1wu9fxJIiqeUU/iN+qzQdf1aQ3Ynvc
BvVbJVEFWpm8Oj3pqrDWoZ35OXMSMZIez75UOavJmg60qHvS/DUVkiqjeZvK40gnhir2JWQIwOo1
lGvdbsP90J5B4WiR8sKDwDBQCaRcu8qHUChyjeb+hK/iB20AE7WX9Tevsej1JNoV7a2gMyQGqExd
DhFqplksrbtgp8w7HYxLFHmeq1iRR0MzzoCWLCeYlW+4ejew31nEmOlxk6Db/zGEqBuWtDIOqA89
RbK9xqwN6h6KU9+vGJQdy5DvbxFKU94NnNqBsjHDiZIHV4T/8wrOJqeBulpDqL4uFxitiiLviLBt
+t8veJ66f+x6Yj8qnxn1Ra3MeM6/+EEcpKA8oxI2ria/8ehm82R/yJy9lA6qtzc2E/kkaRUkRYkP
XmGTyj7yoer0lArqk/cS7t/7hqQiSKzFqcghC2wKP3MsnPRM8yZjIu79AvnbZ9aUWkZY+sxlY2ZQ
/jfstey17K8XHhEgBIzE5+xsBx2ZihUeg8dm9ZOss9WtNYj9rLWG31VbGu5EC+YtOVr0wPtHKfRj
DuWWk9i0v+NQXQgCzs9aWgki1hHJN+X2H+DVhUE2NmlnJlTt9cCvMxG/7P1/rzuCavPKJqHXWB8o
xdzyRDi6nYKgmkpgrhTWTM2qiky8ZydlNXdK7HU4CCWpM06yb46rElKkj0IS/knGmW760jPoVolT
GKlv0JptYb0tzARAmv1TfXJhsX6rrEDTFifToHXUbxvngsX3+/kwtncC85ugXMRzrng5nrOcOpHF
CBMkuFGBhtxtXAWHwNL6pnyItkwfQvohDpHB2uGLd92lVB8JgK2w2O39IP5kNCsrQcmi+mq6smdC
pkbvxPwRA/zDcWkisSIwgWz2SWl7mKj1D6lVyewVM7v3hUJ2iuV93+s+BNx050CnjLe8t7hobrYg
Xa46twAcrn3KD10BmaMUYJ5y+veqWSeCHyLJ1rDuM7IsO3zi0TaHRDk6RSfqQUYHQy6FDgg2QcH3
+joJ5VhXLhCSYAYI/NyRaHySAsUM82yVBzKJ5ZGRLpPaonJJSfxMB06vA5N7v4sCVpqDWfJkMfqA
f53+vy6lhLqHgVk70jESnLwdWetfRM40v6s4iPlYchZI40DO5q7pP6Ol6QkiAXlaDtZcBolCOZ1m
nhzWP708rlfvc0h7mxl56mvaYryijxX7NBayMZZIElf3trkUTTeM9wYHZ5YS0pBgP9N9B2fUsgS8
4GiawxVqXjPjrhU7msiOyrnvdKhcf7qXsNRSFtrO/jrD8e57+BHZu+9DucNNejvpHUjxGdpTZlQl
PtZXpmpcmGlqYtztZnk5Z4C27vx2YLz4LQke1ZAx0z1gtM/vLuk9swu5kiSh8kyVicoFczQ1bPz6
I0kOk8O1C54HQFt4Z3nr7XL1tooMWggU1Vzc0NW1u2B2GSbd3qUZCsJ7l+PhIUjnWS5b6wcaRUfi
PFby8aUnNUn4p/RSSAzhT1L5lbrn+PBSzLSKIXExfSkpk5kO+WHC8Pt1LLDwTm9nlkuuoUN1lH+k
lRwVf454TM3Zd2Z17bAvdnhjTulFOMLlMpHMI8Yu11v64JgZv2Ucy32nKGj6EBIH2GNQWQXsVBOO
KSCEWxwejfBk2FYz5Z55zy7f8Q++vAHkitpmYSY3tj7gGMpShbrRRSGf1qF/HyFnTi5zyaPzadEK
pyMfSk3GDHxQB88yj3/ziM1q+A25um5ZsP2FNjvfCFgcRnptPYQqrjB6YMzB5l0LmXqTpwEktJab
/Fvgul6m75e9Ey9BmGFK1fLdb84kswEm8vc6EDhL02Al4TxqKXOQyJ2dUeOwRPNplzminn3Ovb5h
qU1o3n9FgiPoVvB+LFza2402Pa+1LUSU/CDoF3XuHA75YzHsQxSBlMOgHyNlAJkNGeppScHFETGw
DDFa/fIP/6ER5UP5AuD/jscHkE3bqQ8GD1MYew1takL5AeK8mppoRBCR64z9i/4CSS227Q0gRbR+
OjMqRd2fhKJY0TcJVFHLPIydIwq5Kfw0kxN1a0cYtoyE/RA1rKHA9HgWwxtZWt9qEKnyV/znWbwI
mmm8a0GYS2PB3YW1ndH85ka29HD7abIvxYQv5YPgm4tGThR8YN/lB9GZqKGeLNJyaq5pbArklYJH
Smd6FLQjj2DZkBfxxoaBqtXX9CIvYz8cTYJ3eBwZl6XMEii+j0kQD/a4jNhATEKyeQvqDQoVIC0H
RgqSbQ/Be+Ocjoim26DQ47qsjclnEx0Iy+y00PDGmGz4I1EHcaWUEsevfOPv1Bou0gKYWlm3ldeq
dBcPuPSmHZlJP5Kla3Hg1KqvZUnfza1orVFa6QWTzWFl1VYT90HpobHGRHKZ5dO28jexUrgl87Zp
oN2m1p6rTSbzR4eQjBsNY0Pt43sPKFdNZCDjVZDn4zYS5Ls+jNQwUHqnprxEpVzwS8yzULIsVVbv
LhIxzNoR+aAYOD4aiBgA/c3wUSSnKJ3i5/JvM6PAa1umMvH+bc4c5qNsuLgnIuXhZlDpKUvmRZAi
7XfTg7+Y1vu22mSc1wQRKRzYdMKwVvwcfSQdXLOcknfUUGPGmw1wOvzOMvZROtvyLHLHlzq5zkKk
lvvIP3XHaVyFdEvoE2TymX4Xuj4MOBzx/++1DpTyMRPJFGIySD1te2jCmtdZb7lJb/GBKLOiL1t8
Ynz7P1SGswqWht4eKI53QUS2WhakSsuIuyv6mB0dSxYk8Vvf2T8Y5E2Af42sM23bpsgRdhunT7qt
KvFmIGRKGHUh31PxdRrdPn33DZg+1WQFmnXcILeOvYQLpoVRtxaFvt4i9jVzhYEbRUEcrnlFoq3w
AfCkE0BUFJ+lkN+UZAgGNVzsvktfaTZRcPorchEmOfJf8s9HI/n1L2pE8xKCbPfYHr4zJEkSPr6P
2PJhgsgGnyoLbT11mdIcl8fgGPGv89HdgkjnJcpc8ZcP3bIkliTXIETgZUrJFHsM0WwiwRYTtkas
NCJ0Dw2Z9gJF9R9HjItx3hf2I7IN7570e2Xkd4aASYkfGmBEGdW22fHN5HFbgcV4T51DDwCJmWc9
mUDyBGWOB1TUtly9toOrJJwCya6YrB/tlDT2eLou7pJW0Y0A6jA0vG0MGk/Zt8BktptWvKijEFik
A6VoKAZZmv8kwX1zMJAcNI3bWiImQfDF9V8Vka2TJhX/HdQ4+eFQSlLDytxsrZ7laEVB5rl7PKAz
w7Bm1V93ncJ1E5PAikpdJ3ZXgiy5+oqTvoVnVyo9rGziq8XLYN8S3WRRElQMSqyVHLvyVOGUz8z0
nlZUn/6JiOpqUbpgxAiXbx4kTpQquP4a8XZw5arjWxRX0GsvboaGkfmE/hc3DboVQaoagioeO78n
EkYJJpMDvTUgjgFrYgNk+f4OqkJWKAPhFCZiHcGe+jJC+vL4+LYKeBln0sP4GeyVnQlKXJFppIMB
T0lgO7WCqeIQ6Ex+pFALUvkQIMm4VpJ1GLcmAw/ScKLVuu6cD4IIFi6YIWPncpGyc0G2ztbud1EE
lELUFZkGTyaekwUAa3BIExShbHJKMdjCyhOtE4RU4EWiZ9fxkzuus8yS5RrU3BLTiF1KAyNf/xms
TTHq6/K8UizA+82n4o2XNcYq8gR1ZjFwVaeaKVIonnPN/xdjpB52Zl54hG8wxGi1nS0wLox0ysKR
A1XgWYNqWvrg/EHTZPtA53gEoCSAfGQ7sCGJOVmFyCaeOg5sxBrH4sUUEecObXJ/C37l2Hfwj9b8
COU9WJ70bbXiHsod5AiwPa3vTKzOpOJYGVl39t2fn3iwwydloImZBJwEYDIbnrT+X8Zki44RxLLU
nnlpHu1y3xX4nmUgrvLWKUU0bQw4KT5tB8fzJu2grlqrO/TNKdf++CXdg/g/XRmr4sAfiR+AJU99
14omRfqTvyZDyCr2i5K5woDI6BHXPCmfqDFFP0mehKVaHn/TdcsZDmd0oNG0JDjE9BYfQ4GAC17u
itgBE34mXTX3tGD4xR8H8WM61tIRxo8eVXhmdJHouh+g2nJBaBIYpR2is24HJQQlYXtVLSwXBuNJ
xtcty6q8Mx6xK5MbSEGDTK4JpvMeXriWq+lnGnY1qQWtl7+nu5/GRLdAAQMNO7IPMZBqYB81MQBO
EqmM39KrEJ0rwZyQvuhuvw6JAIeADuko8+dBzO1yyAxnSZTSR1AiljNddlUUmoSRPRnweM+ObbhD
WUybjtikxgz+kBij7X2Dv3s4u8xGvLsZGC2ziFEfFUGsqDF/VAxJv4tRYzNjMqDfQ6C7zh/Yioty
xpOqPSRMZBSrqbzabakLMQMC0sp4HU9NZD3nfY0z6hpk/g3Efkr+yb8VWDRCW7IiodTEqBujFdEP
V817UQ1W8u521RJMJxa+Nk2yj0Xu3p3vtFKefbNn6tX3fzBIe7mWNFZcgbEhO9iQJHTJFeCYBym/
6XclkiLoAx0tkiKF5Hs3lIIEYn2V7AB7ET9SX+mpMmIR6r/oiEpQIzlWD99m/LLvapYygXZ1FM8g
cih4FQ2OWhlu1uimSS0eWa3lhzufTT9S/QQ24STCO0H3a/5EEFfcgeUPJjbgoePpU+UWXucj1LYw
T9juVCPb2xEKnrApQfFA/YmE6xwbutF7RNlO4jFW+5GqUfl1kc+u8AvCEOiQxx8JsoltK3jY4sK5
yyijxth/SL9oKCukHDsDkCTqj6+1Gg/bCkO5NJgpsrtqXoRB1CMiZbeHl2aEQo+K0hoq/tIvOzCp
4joeITujJyV+FJpu+WRjS84ppgVVfEfoAXmwqS9R8iFIC/RvOUUonK9IM7pKJ+Y4rf79Bc+kOPM/
3z+fjGXOPql+YlFWykilMR4wiiSYav27hQqI75Cv+P37jDXYB92UNtzhf4RQJGKVdSNEmXBs0/VP
yXebVMjsGvG/yTujP5f6cCpzcqIdG4BWmcPZisXJFte92a3ayd1viumrgZcYaa5D3U/LZ2lUa4qh
7TFHq7u1myezBtkHeW05D/kjaNEaWvJr5KyhNYSuwGKmuh/HBanZasINA1tRXQckw71+b27FnCD8
fSRz0rFKxavrwzhemNnc6j5NJeSNUyvzNt2/QeLiLU16pcR33NCrnTsC8LJc1JMs6OHPsz7JQ0PQ
gwoo2Yo4hEAIhZy5P4NfbvyGrgldwSRrpvBgGStLCQFuwOiFJugjyplrP4SVwDnVFzUlozO1xGiD
hUOrQMv9ST9vyi13xY0+RvlBKg+Q/bx3HzsUWV4E8k9ROgDnf/d4VCExt/sV9rmIK+9a6tN7QFkd
I5izQLsNvQATqzbft142Lx6Gnf/LeJ00k9J0FIEABI2GoZyZxhi/eCtsTCGLiKBKLgqXSUesmGUz
zZnQi/WpGYMGUvSMWW5tMtWSxq8Iomq8PAmu2SM4hsOBfmMi/7g65u215RbGIaS9F66P6KHOTE1o
8YAR17Pz46HaNbDDr4RqTgC37hJaep/T3Kop9WbEuHhirHa9V1bz5cGESXwXZilSYWo/ry/JCeBG
12lKrtairXAThAZFVoCA+PUHhNdHw2UA2ynkQtZPMpHp0J7memFNhPEQlKAAhkzPc/lo98ax//yn
cUbdMmDh1119GNzvOFOLYY4Uenxeta3sWZ9/NjI49SIGag/XdVl1nbJYfNec/kOGL4/jukBhNuMP
/Bg+jPZyLi3rRmboBHC5ibjtcoDMYd1c4FIOW+azCvY2ohkgTl+sRioYTkRVAD4HjFeXSVMw1z3x
NZNYwGBymk2bYQEjbeUIubKsPFHQFzyO8y83A/WnKLzog6NY5E8nhnIc6yMTpoqBfrPU5o4vC04b
D9LJJdrYGKgDdCMuuOuVrl0UXtSkE9cth4dNiSi65GPpvU0zhy4Yg9IV1sq9Bq5kg2vZqcZJWQUi
rzoi5L9QicMykoYfQb7mKfJlzNKRfp0BW9e084XwLYoor9J2n1vJ1Tiyo4hKdqC7CDwnA8cqagiP
B2LNVUGK82Lc91YorUIQBh+7jkvri0Pwlg9xlOnfoK9/evOpm11YUI2vPpNNZaOi76Pf//8aLqBA
DJqgItyH6xHhPGi/g4Jva02aLeKzlo9LhZ/qoKVy84e9UdSGPfGw2w+odPLFNKchNCuOk/uTa8dV
CW4K54G32H/jU2g2WxTKrkE32Rkr9KQZv13H/YGnegKHknmeXMAo8JxMqr8P3zBs6BB/2Ujdfz/t
1+MTBDo7ijLS1UEsg3hq08q8MZ8lTi6DaJwC4mUn9y11GdZW9h8mZrIxffWhw5AbkLeTcnJ89mT9
f6yo0uoHCzay6gvF588cZnmZgXBV/MfCV2MiAN6FVZSLmf1f6hHvBsWZamjMtshindRBdu08SCGI
qI3ZGgTdiIHDohZjNb/f3AlbluZVpipqnYYxJed3qCitioImWsC153AV2iKmIzbhI84dOYs+XeqC
LPrMTUV/XqaPMVomSyAsIKaHNaE2uJW1NxgPhDS30C6+YHiPcMxt9BGjhjtx2nyPy4BKsAX7Nzo/
x4qbYlkahgnA+dpAEUStYNbq4EgZpJEtLnV7modo0YC0RCX4P85ulyrCiOJ0xabye1D5Sa8Dqxst
IL0bXMweft6SbDKFRwnoJM25Uobn2zou1WRpC0dlLGF1VK/vn8NL9wcfKfBOlRYxflRZigOd5yFq
2+/s3Oxy5cLpaQ1tixWTwHN0tyh/OyinMW8ZKRAqOB7yb5+hOvkR4NphdAaIxrCFG6b9LWJ/X2rg
zYU+369DPrRGbY3KSyjAydi/1+O84g6lEe2ajCw07Ieqqqrk8CNKcM8edg+4v45r7WYzQVzrt92c
EA60zgE4LCtoWJ4xJwxsW64RP3hT1fZpF+39V7K3DvPQ0XJumKwcbAFInQjEFYlkiMORS3gIxScY
Hmi1khA89ecOB4CLGIotaVoTBeSd8vfemZGgxNopgd9eRVL0hBkOUSrnpoBnWGu7Au1Ld0UHeQdF
X0FSa24a4lt39iCsBGPDuOT8xQrxigIt4PTq6MJ+XQky3airH2PX2dg34OdAl8JmS/rv5k/Yie1M
lbBvQC/Gn1gW8ZjGXqt9lKSE3WGowmZ9J3B2EwfkTtwIxE3fBMI0txJR0A1z0oDcT6SUN8XumgZD
wqWeMs1VIaRon1FGrSUV5SR2cfUVCfHIj9/Rmt0LnCbaS27X48LU6uqwpvZkYyqM4/kOiUKai2nb
CxWA+bQ/Ez13+RL5wruU/RO9VDFQsf36zrBNEGi9YzkFc2rzK1iMsPohoNc9ukezly7sbfZaERIB
noBm63Fa0dD32a+2yhr1AQVZaWj4HUIyWAaQlibNMgvz8GBcW/tSPAYsg1cJLxbcNNjypQR8LlZw
nrWfkSkMPcWQYvpyRG2KD6HtDMOhan9cIf6bNg5KTlnqVZpk047kFrAu1brh8pZBtbKKHnSqUJhR
YYpfrsjK7c866PSUfDrAKii1AEqdVO/wvB79BLaylHSQDzHOHtP/AH2lTopr1bqpkd8f/3dWaxdo
6g4M6/fF5jzD23eO+hfPccQvGINhyaiKO1w5s5F6SEJlO9IEay//4xWe73HHAvrwCiQbb88HY5LV
v65v7G/6Pb+II+yGRTgWa5hEPVOw//7Rnek8BXJYeKKfNjwDyW5xh0lI4EIa65VWCEGxiNn2vr8J
YCtSLdb/RpvjKiVh9fIVU+0Z1JcveAGwaFk4XiC5sK/89ZuKTQ9oGsdL5EAln0Y+ZslqmKuREqF3
2mICBrenVejZxCcEgazUs20IKw4y0IhWqVK7tlyf2uG/3ic/bvfATph0wFZIKvkTgEppFNXd3WF+
7g8CfV4Db+KMOms6FexX+WEUXQzzspYx8sOugjSvohpgdnx5UW74jJDaJ4hPJgf7qNdmsSfe4JPK
+1cIWal0z6JVtKNBxfieU46D9SLFXALy9lRm93QfsPNQGVUobBDq1flCb4+tdZl7fqvYjAINyh7k
EZYiMPFB5SG/4JG0+93ss7IGbE+NVDp5SqfMyUM6BaDHpKIUpwsCCglfcUqmyUxJ+7xAZckX/v8r
NABfyGPX3TwXXsLXd1y1AN5hE43eprTfnNtUbUxKzSlDuDIyvW84NExmXDuU6kMd6MPn5uCwFYQY
5MT5pxL95IPnVuDxGw5RYQ6LsiJCeJFrN1E8F51j84w6J3GCumC/X4XCR5GTvs+4HuxB+faW+vMF
albGpmY+nhrMwd344CTEZEtNSEqDTAG59bfnv5UqghocdDmz/ansjW7QVUsc+RSrjfuzN4N1X+c7
pmGG09hA4ONbudMt1OlarHFUWfsewSgSNQFH+ZS29OJCfJRMCd4QFIHQVc8jqs4xDxoFO19T2R+F
UvVv3GMMRttB2ur4hY91j3gj+3rENh8trhrTDbqHMR6g9iecHERJOmHWIR5S4L0HdsxWWMQ26x8A
oP6tXJI6ngn+Np30BoE9bi/Zxb8B4UEYtm8pN/XtK1nu06lRi3nCRxf2CPEyX+/Aj61md+te0i59
U5yoFk0a6fFnEuOjOul/e1TE3FxKNYIDoi/zjA7x314ZWj/XL8MDVu/2FH+1bLplpR9KqMAAF1MM
gQzDE8jzqxsfHHipZ/lPYD2MKAKCGA+wwhexNz1P5SrkPDGr2vgzuN24Nqd7uxy6iXL9GHHrLNx9
Jz3SdT6ZtfbQYIGiDyvdmVD5M9G6fz53aAF0dxzSyaoev7LxgtxLXdCIvRpIdqHnSbe/lygyZp7Z
ufdP7Ax86OzpMvhXHZFRiX3KKDnZXoqiPS0DgzZJJU7MkWUKv0cLwHcJYYs1JH5pE2al2Aw6dMnv
D1ziC6wxOgpubxuG3VgkndMmHLeSwPyVgEXHgAE5Rl7NF/7kfayaq/PJLegc2b6vx36713QL3H7R
9Vsa309bTm5jQQ6sOxxj9OxIl6+6MaYb2coYzj6kc6WcLkDu9kxGb+QuWK3fiX7AYWBn3uQ4C2Tt
tzzum7olc0bvi9vPLiktCAyNz1D4B8/JhCfE9mYdrEMnqpoZehRPn4JgCzrQQFgZPpm/tWQ04sIv
pW+Otacm0z1AZH9Fk/lHZK8VdO5x51MFoJCmUzTffkQ2XLRIxmAdtQ3YKkhS3iXIg6Qw2owpKTL8
KpgcKdr3kR2GVg4QQq0ZKNVW2NUger7UvmPm7TIcs9uwpreq3R5t/PnWhvEuJ6J2TRqbWIeEgZ5b
ghrp3LNuO7eOvgAzLws2XsNRPBcA9/tk7CSDRad3LeFIX1G0J18zVaDSRd/88+cFXhla2+G0E7YI
5X1nGWAcU2ZIBRVaBUlzzfSU9Z/422ih0uqTaAE1ZsTLOaumhqKLV2p1mlYN9chRAH1Jgu9PI454
fYqoKFW6+te8mPh4/zMd17Tj+3W9xPJbnsezNN2zhWe3X0n+6aUmz74CUJKrcE+cVcvG1xWEJ2wG
mgGo82RFCgmq29HyfqeJ+3Dc9ENMURBm9bfEnw5JOW8KRAUvnchc9OomyvAyLv/7LbPlxtUCzenT
AhsTou2jFv8Cs3BTb9XZcziEWYd7008pWJlbzWFGaXeB7WtiOionC11dgLzn/bfSZ487qxpeQTQN
3rfz5op8r9i2BTpepBBMZlGftfhAJTsh/Ba1+Lna7wGvtJ8a31QzGXUUpxXpwmo1V3on50ucpM//
Q+F1biV5I9rocKH9PHrl24V+zEnxn3LDCqAOc+k/1Y1Wv3qD4WtENf9lm9bXBesxBscye3IzUf5+
Jdsl+Ds9NuZHJujEABPaXRleOTbmqFRZvMyQT38YKybmA1oMadYfIL4KFMqWy3ll/8bYTFG3wlqb
vUtsFXuY7P7JO8ANaweIOg9y7COIQegjxDR8xkIO49N313UT/ejUJFgreEKLQsWpiLDVsX3zOpGr
E2hwC+ea2zhtQSa1Y1x/FFooMIqs1dWRUVw5u+3ssi/71R28jML55WlyN3/PW70yu+5MDyk3Cb6l
HKHaHDX5C84oHNKNGS6xHlkaAxwLIEqlS4vrhfVckhm9jpFu6jcq5ZZI/E89a+7MHWZZEi8BPmkC
WOyJd659Q0QCebVOBXNgqvITfb9PDH7DaflG5yhO2wTUn8ZX8vNKPiyePP6hlCxO3w0prxRXZg9x
vSITz006/qnbK4VbouHyO7wnowul32U3xzIRXl2A55OblOI4I48UkcyLsb1RVkbMNEq1ZzZQS1g6
z7zGJIAh28tDeSJmoO8aQGJczhqNkISGVNfIFnyfKjSsgiuUasJM4/MaGUitObTrsRVRLlZ2BcXt
NHVuJ8zglnKjeWHBtDMFf9RhFVeKj4yLuh2a0D2O4JYh4a5fiw1CXMLAQV8wsby808+fVVTa4CkS
ojNmom45o3YDxjMoffNhwrfky/nSbXOS+xeDdaoUWx2Vastz1LcN257wbuwjeQAfRoeMOF0NkmFg
5Dqkp4O0Vz3cdkdPwip+eAQzcXi4AJ58745mCz1uE+ctQw0OQYd4d8HEAKaxbhlEsmn69dhZHhMP
h8RYn+XHAD8fRAF0qnFiAzTgbzkhEu0KwVPEl3mCKlMeDsPkAqYfAHOqosmbuApjI+Gh0aZco7NA
0GMe3rhQ2ULkCKodKTxtLfntUsvKymTbPdXaPxinTVgf0Gmj48txc++pc1K2zWUQQG5ZFdI2bAXr
MtybCgh/NNoaG3r9oBFCnkh//blxKA0PnMV4vbfNdWHT+4l3IfhijCPVooStIvvIv0awrVXPdrxa
idKGP9okVIPPTE0O/IO34Q8uF1cgWcOOHlg3Id6ZUt10X/k8ffYl0IfLDSUvWb0s+kKgeEeA/4Z2
5XHTDyc1tPd1Nvgd0KmhhYN/NsqBsFT7HRsDSYe4LBQ/Blk6y61KR1bVi/uP5DQ5dqlnXDfhPOcw
9/YJ19zzZm45+TzuMAdAVTkwqzMJ1kMvRpG9DeZEFuFyk1Lr5Eougnzbwqial+sIsfihdOUG+Az1
9HUIHL+nYmrjIB2FKiZNy4BTpJrnBS7sjLlFDekIONmu6H1s/M8xdgOaQZqoyyKzikJp+gRmKx2S
L3kSLO3x2y6RYAH2H7Rg1FaumPeXMu8YEnCT6JaEfrhn5NoEMkBO/nzsW60dx3CteFXbcfav//oT
WOl2nOcu0tXeFaJL2Jz1x/26zBedPtzz+PwS27sBwsHOrHj5JW6XPbBbws7B1UkFZ1xssodRt2AV
s36cNIan+7HIxY6c7ypv98q+QNmc4Ac9bg5vmgKNcAZ3CDVSCN1cOYWIMKONZ5d22V9/dYPeanHa
8Lpi5oo9X1QhgEUFUr+tauR5mYf5pReOrfiR472oE1vuYUbgmJ+QULL6Xdv3uvN6khatiDNNe7Xx
olg19GUO4s4ZIviTBFy44yIWXMgGQ0HSbNO4VC59r0tpgsDwmO3anFt/5Y12v8+/mSUIQzjKK3Om
Z7nmkL6E0rc4XWTsw5SBeyBPz10HA3i6RSUtQInF3wxr1F+wyL3djbNMHgsKnB6wbWSrykf8Eg9k
M3p6QCWTVAATGld/d0l9ftRlGewN3uIn+KdyRX7RFgVwmZWkIUF5FXcuVCOnFIV0xpjr5mBa8Ybu
zq/OyiBAnjOEB1OhZoA69KSv9FfnFSqHu444gCq+ZjfNUy4rOf9jzb2O3RMEZtiOXh9vdu955sVG
zjs5rYcaXol9gpieN48DpXFzyAtkoY3TY5cMqN7L3NXanfX9+1GIFd77ltcBZ54cRtCMIBcE+coz
coVdmWYTRfPrDq237hhU6H3/WiR3uLSTICoYTKJlZ1Dmv4GzXxYFFFUi96NRy2qLjYnPs0jW1Ewp
UwdM/kjcm3wB3vaUX/+Nvj95/JtW1//JOjQelc0ai+kvxLGaM0BCRoFsit9e+KjLzof8ZMIyw/yb
FglGOg/FauUAsGXi6kM6UC1OEZ5d+iQcj5z2ETf3e8lYYzlvowInvkRfpt0pmY0E3axTOHKi+ZbP
hG46gA8wVm2FPh5DEzgYWFP2Qt4CngdjaYiF5lq2WNwpLNXfWchgWcxFJ2Dw+yUxzAEHcojDKtxf
N3U9xxQLSTlVfZwocQKQeKnTR8aCYRKN7KN9oeDt+n+WBnY1/xiAY2o6Ngibt7oxHIIM0oxVAnNS
iPIdw3F6kiTuB+3SOXlcTxNSfI4beTw2iFyQt1ToYBsWqTOqd3qWLPwtNOlzHUPw9X17xm96E0CE
Ok8tSbau6CrTi99o5IOocMYAEPU0vvgNGwiLU/vxcuxeSRfp+KFBkmXn0XJxzqxtXFEng+icMOwR
TD2nWvdeZ0Ao4Efwrbe5NRR+PxskMOH3l+B+IHncoSWt7Eol6DWkAZNkv8l9uZj55oEWsloDtxzE
ajczLccQFPv7ST2FCz9MbvcRt2ZzKLJgXKauPulPIzXNRHU4Z+/IxqL0ql3E0F1LUD83d0rvl2vO
clJHOvue0hEGfSeMURGNdCOAbOXld49deC6NNzFNY1h39wfUcDzMVDGeBEghl8UuD0Mw5B2LdDPy
kzAL4zIZEK0cRtGDUxEClh16panMAyO503jnSINojZ17WVW1jJsYB6QjVuQdXFH1RNkuB7nkj1NW
iFQs1B6eqlh4fmcdFGGVmYyyBrU5eyelPCqL0EGUeDclDY7pKhpGU+1Yy8ZOZAzYvYo2BmlTVJ6r
5W5T1n+u+7ZJndXfSS1RatyqvzaJzQqf2o6WsIgcXiJJogRTMDKi8nI9ByEaXYCAoSeRRd1GdGrX
d1aQNcquIGhBcFHoxEi4JiCgCom6hRaZH+zxNdCwxjdLX+FFY18mCqWrxQ16MC1Z2+zhI0JT4HZQ
P5Win0Fe2PvgwUuMHwwB19R6voKV4Z+woOy5cynmewZyXA3AjlS6aBqcfhtAT0hIaiE57O6HtALs
YBONffHnvtbPKVWxGErCLuHpAyIonqecQ7njXWSUGhnigxeSvMIFM8buKCOZkQ+4N5N9HIYeozUe
TOqQ16ObO77wTqgyJMdsDKmLcUdJuH9WSo1x339eLeIBS10cocVGt7tQadteUhKvNVl5J5QvGg3z
uG5xc0ACLE0emxD1W+CevQXTZ99uX6ZFmxHYq8A9H5jKEnUtchxS9HiFYygbXmlsAm0HdIh7fNMX
y4TdhLUp9Tkos2WHMonZWxg/AXSm7HuzRUchqexmi1i3BGFwwp7zfXU0bPhx+jKivQnm9gsYqL5l
+OuFJ+6/+qZLq9bLVVQMqGoPJwJLb39DGbj9GPmiIMgXUMKzm0lD84xlUl8k+uAfCp2p5ptslYFD
RPrpj9nAMiFnnLmHZ6yMzzUhqmafzHunyR7TqG0k7aDs/WRjIPuQ35Gn5eHOEIovgypAimkS41kE
aJmTOwk9nH+67cjnruh0EviafkRfhOnIxJ20oj0e7g3QBROZRp5CcdmWXxvu1KDkhtuaaVe4WL1n
K8VRuQJA4LkJCBCBAKuo90OKF9cO3XUDGjXY8wYHabhqvOhvcXJSQDGvC3dr7pCb0itAQgrZy46C
u1+3iY6wrv+y7zn5LFhRsnq7+Z2l8SYsGLkNTkt0LAXxd/C8Vl7shDcMFeKP/CnuLWS0DkTjuscj
twq7BNDgM1wAMxiqA+7mNxmYP52rtYzRC4Hy0jhHc2k/+nZtdydWKKJB8FnKQzKS4w68VcHUoUsT
WsnquccICxMNOQJhtsDWjy7cJ7PsvrM8p3WZ56o8D+y9ln0dTP/3pTKyFY6N72t2fTcnieQ5GGdG
mJlYAaiwX7shY7bS+u9vs+RDyZTjz2zPHFnzyPY7rqrtsQOf3TC8bxcxsSRTj49K0f0SKT3cXfCk
VgolcbxWTwIovS0LR10zQEMbXv2BIbgEDz9FB18y7EbuJ9HxmDqHuuFC7A3frSvX+a9hqjkHpooM
pE5oi+y5VBMDRhso1fVb9A/CnAMAOvPt5pRGmxggdcTppFfuEv4Iwuimm22oXrfSo5sIZoiv41E7
K0kRr0Rv8ZXytxb60vcftOZcT2GS4nnvrrnJPivvU00MgrsfF2kdxt1+N6HGWOE1V7dU9q+qxsq9
8pbkyzQRpkcZ6SmQswrCkqxzWtBRsFOkDEoUeTx2iMNF+wac7oIRB1U8IILNBoRYY5fvLZvpolOX
NQTryhclLLdbPc9bHDpVPT3pCaDVXOYDbJOI4BJa8EYf2JCTiPbw/+SmBZl3aoWZKgCQ6YfiVzhm
yQ7JWMeOmU3doN8Er3V2dZXAQXQwZYNvgxT4xH05L/VkvzUtIdWxCYkV8IpW/aZLo2UKH6x9hilV
xcz+05twbai/nN3NbB0uG5qK4FWnqz9tpxkWTQGS6yr3dfaPwIYVBLmM0I44ZMq6mkMgzI5syT/L
X3ZG1ScLUNNtkUgUJVrcuvgz+ccQXh5xREoXDN/jcfZGZ+0lHh2f2GvGm0kEvBoqKITjqD+jGKj5
O5wuo9vGYW5ZoWmTparppGZluyPjNgk9yZ1gHxZeb66GwJ+QtP1eN9q5I3hMcG5HbVOEfT5QH0ZL
ZczbmVkwCstt7iU6hSsS088zD0MewMGLBBcl2/QsZUV2n8mkMgcgp6XoZlXnQRD9zgvfjb0ac5x1
YE02kgV2z2gSI+PgZmLzth+KQlakMGTGzmG/T0zAwDMlMJVsCZR6faSmYbY96y4Ou42HR7QnlGF8
2WxAxBF/AD/7ePRxEseXzPrhuoL7p+KdBxWWtQ9Q+BPAXktWxBR7WiBHCpl1pKu7PHLANxNaP57A
pkkWpRGj+rLnDrr0jhIQGaqhT/TX+i8JFxoSfOaxSP8TpjkJ0TGjlfl5YIQ6mcZlHVn1RtrvJRZ+
hM8WEZwGe+QX99tn0d/3It3OfHvD1SK0deRZMMLx5JUcyZ+IMw43q75zjvCFYkGZM+h3svrHhJ6p
3vYXDRyVuptjrnN7ubMoaky0B2ThuFcTrlIu7tCL33tc6YI2lUo+d22+FBGMj1fIVjfzMOpvT9Ne
H97lu/7eyar3INarmilIgSnNlyoHDSLDFtCaQAMlAzGGToZ3tKgYXs5ablHX30oWKgzNSLcTM7VH
lAv26356aZmx66OKqkdzoDZuK4vl/p4lUjPa6VWFUcvZiGJr12gKgbqJ7DfHIe4InHCY3SZ4RuWQ
1rDBHe6Z41COE14N0/ATnGwhfWoUS3jUW3YLP7wbgX+WM2F28bnYogrsJ75fC52tutVKrogC+i8p
bPlFtvLojcZ8m1awmXsltIoSSATOsUs6yRpOFVACuX4fo1mSAQkFoUqvbdnqxw4Ez27rD0o56aqX
zhmsmAoc4opdy43CNDEIT7NrCk0hGwpIYR9BgF2Z1FaRRajIt/zEOQzSBWt3+dBNGy9a8ecVG3W6
YiWO/J81Y0phuEJnCw399dJ0A0hm68FFtVxArsXD/kwCogwUzRoxJRsfmUVE6X8Y6ZmkX6EXhuhO
8BlLwqYKAE06/37ntVcjIV/u3f/5T/PGfkSr6IQZ5Tb2IFyNla/hPI0eJmbCPfAzSvKIeVRDkGOh
/39MDDuFmib4whEZG/gNTqlbekmk10gyE6inDbpiV3wcyqCFDqHnhMToT+ySczARvz9XFzK2Fl9X
7K2qrfDsyCdOKar1/0QBS1QT8dHh0QmMnNGQ5gVSj9JEfj5JweaKK9lk+36Ws36S9Y9oRox/oOtr
OIyi+ar/feAiGDYF4ZryB9PCF4Vsdksem/wsDQSNLF6sU8ndh9AxwXWcCYJB6Q3IgHpvqzjvTMDY
dC4xlOf8x0cHRdv577QN+CeltbN5lOBeCwBL/AST37Xr9UCtmyy4yWf92JxgYpcUFQVmu7wFe8jY
Ej8f6q3sY1JnF63VRaOq+uLKp6Qyg0D/r3Pt70ihuIzKhU4GaC+B8qQYrD/TuaJ+52mpE0zU+ZLQ
azjq32CcJJcYcqKjk7qB6FhMWR3/pWzNouHBt2wBLeTuXrX+KEI5/LNIf1l5yWcc16WpLrOhMLGB
oUaMgSRPnS/hpdXkwPvioTy5m1PhE65RBYwRFwYFGlbcc6IMAuzXexULMm/hJSUWXvW+SLslbiQE
uCzHJBMFdx706ybKvNL8Wyr66Ln2uc19GWnqg8dPbQRs51f5vVNU2HclkaPllIlcYligIUaKBDQg
HfKI+NaD62hmRTH1b+SPNFXdJZAf17c5tJUr0otpztcikb7zYHXrEhb8AA+INJk8wseES5SQAFdx
v6Hf/rulNzKDn/zyJTDzkoHn4uP7Kbdn1eCPYnKrXZOswdia7qlsjLenUVfCT7yAfkc2WBgmQSCg
epYMddh+Zx3nwqS6AFno6cqfd+akoAQigg7L07Xti0NkYDXP++xJN67yO3gWEpNPHviSEsTICHzv
P4KVl7+bCn0PP91Gr3sNWRJKLU6ln+2Viqn2Njr8PZtnWN3aWDXt6tfMleqHouhQBmXRJeg5VtYh
F55ylWfCJ06GA4ynk1f0n4yZaoc4JrmjvmXTtcwrTriEU+CQsysQiH0KfkkfwbPS33zoK4puKXUo
/De3YjEyI073ugZ3xGYLFV2t4xuf0sZ9VfMTGNS38ygLdCUkYnURhsduSHlcAj6ZFHHIDWwy8cfD
BtdN/SvIAqIv+/l06uqEjSTg5zl9vPrJfpWvZGLMr66/00skORmP1OFlcsv8FH5VQV91JME1jjDo
9m6bRTOcD2JxiryYOWnWUDumVtzuNlPIif56z3LxYRkw2Sm/MMMJ4Ce9/8r2euOBFvv91wM2Jmqr
osoOKG7aiKeUB/lge/y6YON/Hu18orWsuoq2G2ggF2YlOpqcJ/Lc4CHti656/OqG+SSI1fgDOPJx
cPTTbDl4xz5uJvAQCC9jmkV5ZfncfaROBDQr83IAC/43gxbvXPuWrjnkz8MqBMW9kCb5DInA+hI0
YK0tPcj7WeOSqcXkS41NKNW2AfIoSK/34CMzuzLYjIrj1HQ7iPDq97732COxAX4xgvz8PYhcf8YI
50izibldN8doZSFuAvVmaUHgugVwPyPs9LlqeWbsY2YOm4pe5h0qWSYz04Wwt7hlWxrUb9DVWIaR
Em54XoCUGFlpt4d5WSX+vHPRNqCJrUt1ptvp8v56sTmvSEL12hItkZJ6H5uxND6t45RjL4EanihP
ap1HxnU1A+opLRmquAhL6vPwoxSEfvFwCsKGUi3PGLYX89FV+MHze2Bw7Y11+OVSHzTluXL106M8
MwDSSxVUMG8QKs0nTXSRktHJxxac2TOyIXc4v1aoTOidvDR7eSKyP9TaeAuA/4E7sTUeDXkqk8R6
fcQjFIsSsyvlo24clSMAMap7pYqWME3moObqHTg1fvLuAOHQbwy6tZRHI0RgwkmVRj9lJhZer01f
toO+eXBQy8GCJgBDSqrnvpUmda/y/gVIu30zIv+hvCdkdfHA5qBvwWRuifhuRagRBBAgQWL6cJzy
nJkgfteuyshpyWnIpA3ZyBvSyjViDZ3KiKbe+N3dpYR8vSXMMs0DbTE39QcZszgz8zjjk6zEwMZn
N5r5Mhmwlg2j/6QZl1RJwUn53TYc0rw0pGAuBbqE1gRQNwsek/8W7pM9z92sL1Y3o8aYA4IeYi+h
4M8sJwI+9nFJ+TPfuPKqqC2iqPYeCdLkN/HIloETA99KNmB6PXQBz4sYtcHOiLjFikc+2MkCVNq3
YQYB/+XQS77++lQsqOK2kfBd0qp3TMTfRRlJl9Z8qE7IPrCLRUhq/FOtSxTP8h7Y/zsNAVEcDfr2
Fy5LojoRxcL4etpkaqTGHSOaDuwXTtjjFQSUlVDTPjJeZa5ks3H6Qe+dnb12yQ6Dadj925IXAUNj
t+EOtTAQb/ia1T7UNODTU8XmRaqwGbq2q7MGdj/Y01P5AT0KPAHN7zlPw5TQY1id2Li6w0E8xZiw
DFqVgHMQKlbuo0cRM2F+InyZ92SAqgxaJxqDeLDyTxRZTWjGoM5mieUlb6LhzigGGOUoEGpM7h89
fuuA8USCicLVFY3UvzK+B42scuPEwQOnMH4BYvPKFIjdDsBeVCjRjAKmXxMtI79dk+ZJ1AM09ijZ
akLnmh7JV5CMeIcmeAOdRIr3s8AQpXXmwFd9BSzge0emOpc1ZyQeNOoNiRUE/os+qFxjhhALkogN
319a4hME3EyXPYQMk5u7PDw/euBp3pEQZfoVnEaBiwTzqAGe5n4lSjSfqx+DI06BciVmqBoHqgpu
y1RS0YKtRBZn3+jl+9P6dRiCYOmG3rXZW0hidp0oapNgUzcUSLY99AJtJyQoQvwTjc0R7m62qIgl
fA7fHsCjiGwKMkgeU7cY7wJN/J3bn+eF4EVyw5eRCNBKTtu6hDeDZDSjwbIBSbzZa8+aWg3YQbIp
Ok4y2dTU8PgpZRTe+1mKozQBdckgiSmP6maax50Hrps+q00mGXtuaioScO7Q51/MCXcjSPj48nam
LCHUbyYMyNb8CZKgAsCBhZHbe352BOHaCVmyYfIMkbCrqDB6wvixDVcUAJqASN+1N01OaRdcZnCY
0nNDqlBq2QTqwVIUxZXuKPvkpDX+lne52uInDMxxBClJZ0yH4yimNGBKh6K15YRo2QOBLXzaY8Ko
C9POflQgE79JZpTzUhIVSB+nuAyOXOauUEQIgoAfWlJ8qAIJSmB92zK3JcKtJp58ybLexZEWqIFb
5s4bmmzb22vJWPUfKDHZjdUni9pzMSCIBTvwdNbmpwR6XM6e0L6lYwqWl9gf8nTo5jjhUupHrDiQ
7fRW0o8Pap5rfzOAu1ARJCRb1EytS6eVe5CDrShP2LNnuP1WDDFLGv0lwrp/4iUKEp8z62yPYDpp
rME6ia2/kjqmrH/13Bqgc4UcvkDz6idAMYXJUfeq3ctPEfmrmPvoQXhwW3sT6T8dCcZYW1hYSHDd
vNkoBr1hgz3+W/jOdv9qY5RZjE+cODOAfK7GjDQcGhS3BZgkp1qpSH1xMg55sRl397fWid9gXUhw
wLt7KfHoxQTL2Cr2MXhI3uN43iTberqaYXXDh/OyCiMPKIqNutIZ/PEy7xLIiiDX2bPHmdBuzcnp
k1XCNbS+RG2ZQ48l/uCw1xjWoZNeDfxnBNvrxs2vj88Cq6vaVQDlcHN3sZI796RvaU6SsJOh5Ihd
SKBrD+7fgq/stERs2STUY9tN1U6CeziRdwvO6OrwQBnxOa1RUjgVhKJEFlUL5TNHPKkkvLoWID5Z
vVAWc2DkuE9VVbUsez1RtbpMsZptyrZ5lXgAezgPkJ7BhZaJFIGVv/lN1e9QRD11AXinv5MFhAlv
MNICYxDReXcjrvFaQIe5VTt21T2Aetl3FSaVnSz8jXaT4ZKVUW8sxJm4q3VsqPBwdYtqZaZR/TyS
EU0XdYceYYN+ZSz8wcuSSXkiySmm3THXrv6aDIwnvhM5Zc63KtUUSLaZYbEAt0SlXoYMkkR0ucGW
MZsEMtO5Bf6TFp5AXr1QW2uCFYgpEER9E421fnzFJrhGvARnvMHFuBUJCL+AQiT3oYAu2Ixix7zd
xmc99fYdCpVvmhw9myeTXBtYBXQ5diouNip3Wrg4aRPU+62pNHhAuZ/CrW7+8+mPnS99cWBI5ktO
nD4eA18LTD2+q0iuS8/oUaLhBS66295gJ2weTOpm9q4eH+Rh5X0fO2Lkk8kRnMg+zzfcAXGtVz0t
zdQYndwd7GsxjYtKVpd9SZraAla6siOOwQB69OZWkunza8r3uR/OFKTy4g3aLeArSJ2mtgVZ4now
jojB7K/T1C6rCi4BtwQJtScZ9G28w7dUtRSZXwS1jZJVjS32D1b+qJi3kTcCxCu9TVCCIWot5qMd
S1FhE5rdoGWQuRa+dmlGZLY4wYNAAyEuAuJtH8bRPIUFVEvhWEtPGrYKFqTy79EkjvxiS9oKiDAb
Zan9Dg9mFpjdeFBrkok+zIkj0GyL6Wla51ZDo7KlmrIRpevYDNlOuWcYhNd8BrIlQv3UGgE5HGhS
0w+BL0IhcGtC/KOszWK/kjTbDcunFxWt7NkO0Li2JG6TYJW5BpeEHUsgJIKr0CwQECHJQPo/Sw8o
O4sYabi7zJX8TT6idJQPXWd44KOHeODb417BcdvTqcx7g3ui8pw3VvUyEe7D2sGhPc0E4dbGnSHp
OAO+MKzIqx5g0igt0S3yAYiqqsTZ4DxQiFnrJ6bnnIpfZD2jtjaCixDxhDm+Dg5s9b8rGMYZrxDi
fB1fxzFV2rgRryCOJBP4GPtHf2A0evBJw4yadqJ26IFuuFUIyCSbNf+XKqIbKv1m//xBzjs06E06
OaH/ejBxWJwqryHrmoWHZ6ARqTIA5mREdrPO4cGeIQV0Z2G29P/RPgHuXeur7Dl0zXqYYXgfrO9T
9F1nojN/ZucFeSLbLVR+c3fS83LKKVXplVeMKjJAVafpKrzjn84uRqeUQx2frVGt01iL8m1jgwo5
7M/YC7zXULutiPxceR+EvrHWdFeg1gwHm095YkTJJ2hKrh25eiowTSz+AqL8DgDXrrJ/eAZxkNB8
GTQhEWroF2MUXnAiotHKckso5FgWMLkYLWHInaphQs16erQnKEbQ1OUdPWPdL4wX3YlHpGiRtCrZ
SwNLheNkRuYFCO49Lz7UkV0/topawLV8H8EkZ97Dt2x6QkKG7KvjbKLRE2xvoufMDwonyfdSNhFk
bBdjIrEKhq6CNE4NnRtbSJPbXxzP7qbLXLlPDPiFy06zL0PFfAW9JAF0+L10ogVqSQfMyf6TUrKm
Mei9jTlMuz9J5l53R7Vyyz9RvwexRm5jMgwz2gky054Bege9x5kYqk1OprFJDyhLa5teEa/WsQ5F
830bwWEW9qzuA0A3lwb5BWhFhK3brAdlcvSUPTWPMifDD3wZxWcuzj8/Oh9FInfSdK5cJHiP3/YN
AmBmLNqKBFzyq8lpb2h61j3AUZPw0m/8kwRiWihycrXVnJ9/qaXzV9aEdZBY9LN1vLW8dYIhK0FP
sSXibxZQzb94/ptCKEuzmEDt0NKd+OSlnnWmpZ7NDgyheH4XVdSdi1bvobRNTMTK2GQJhgiPZPo+
Y8fp24TNYSl53eZW1CeA/6twpeBaj7RPklLt5fneQXtIAFQ5L3g0C4p7+S5H0S5yIxs89ytqHM+1
2R4qbHNevMQu1ZnnUaZv5JcC4tcaqepwwUGjbZ3wULNNEZDYzWabf8+T8GxZR3c1mDph43jyGieR
OK0/9bf39MW977zMx/qTQnXRlKsCAQX8n2oSKP/ExHeCoVGQD2aI2/tBexuWMARJrznMpnHUpH+o
jmy6RpsYBc1eRgVPr/2vteo5PI1Jymvh1CScpl11bEHRfLHSbVyHPfK/0qTtoBsIESyRr/4fY1bh
YrmsBlh5+hixKLgnnt4q77GVcj25wAvtpBdZ6jEWvgX7aH4QESf+AV1m3WVPOTrDPgoRzFojUV01
8YVd6ZW0wF20Xwap8kEzr6BGhq82/bTpvjrPMxOczp3yskH+C2rGUoiCDp1J9o3llZi6qWryALVa
YD7dphh8vadMPJdOlMIEqu3e2XXnDuDytoGhcUedXq28UqCixydw4gImLQvHZFNKAe7g9OhZhB6/
NhaWSg9rPKfv5tHLnGpaPfzgRAIK3rn5k4HJpbE1U5RvJ2W2e2rhTrjAZoi/XNVVPY5lHG+luuCR
BZFrVBn2t3iR2Ww9bNoMCCB+/SJ1HUVpTyfrHi9SR4uGmi1m71nzrzZZuJoC6XNNRAO6TvpNHIKa
ZCRQU0HhsPSm2xh5gy93iQo0p8PlcxCiYSXwJxdt+XOehdqfa4jkHFqbounyxXiaOMq2MIFjC5uI
P+w65JI6IWi77sUMiwB5Y3qLPLDlQXLLbfjNpJE4DcIHvkS66JMd0Qn1P75n0UbwcRTq2gjEsd+1
LxBsjc2sUbaenidHEeOfjtg5UM/ItWAO8HScAukupw9nWmA0pVoMeTPXP4QKO3G4HUF5x4pmpLCV
4juvb/kVKP9Eg5M2L8f38dwbt3Id4AlzUMx7a016oJjYgnaD29j6H8LZBaHhn50xHW+nXOjCqtNl
Sb9MK4O1MKmVd3yIQTPVfgKCmgQhtYAlLy50PuW+/D5LPBX19KveBVyVV/UPagpDKf6NFSXkxxZO
ecskyL6+TERwLpBRbd+dTO3z/ZuTnKbt43V1e3aQjYVQWQ6H9DHjIU6vZ3R95Izw7CikWRpnXErv
Z4sdxzlmPcx7Q7+GlCB5+WYfLmuTAhLvrx0L73tympgIOPeCAVTcIqjUCQRKxU47olpRM7+2Yyon
qqfgtStoTCh0onwQOGlFmDwlvkgEL8lDhFmr9DIxj+VdzDy5Lvvz3zwX4VlWt1DbOen0PlDuKGkz
qNr50Dfv+zkHpxPbj/cS/Ilx8gEHOTCjSur5hnqt64/p6MaHkA2t9W4E7Oj7f7Sxoq6Jn98VwhvK
YiK4JGuCmHcsZLWEqTB2iO6SSgSDuKXUxpYh3KfX2z654iqWwXw5pZWHC1LgOQR7OgSaTKnZ35jY
o9kVZhO0BV0yHLtC3w3zwUyEFAEibGqOepswrYCe/IOn7PC6Buwi0aQiDsQ1qz5/Vk1BoX3dWun5
kncsQmJWJai4zwoeleIziCD6kYfrfO6dHJGhPOQI95lCk+ZtBiFrlCIG1+ufeJ5nmv4ixMoTlOVb
8jF3meCA21ZnC0Fi0B/EO7mYTz58Z1pn37aTi91+bsLmYearX21JRFLXzD+6+QMQrfxBEcvplrOn
/0oy+0FzXz2S/vltSn1MNRbEyVOch2ealVSenlwMPzAp5gAn6R0cJ7Piqinb0xfd31RyiyQQhJP2
NtraBUJEfTevrOMB7q1npS5zfbk2vR5Pm3hEdAzjMybE5sdcYNlwED75Jg1OIC6wMwrRDIMCxKe6
caPTBN/1t8cVlYB0kjb1pwXO3B0PlEEQVhv75UihPem2+75upGufVPUUhwcMlU4a0ex7UM8hcDVU
5RFMJMwOdu2gFB+tz1wVSU9JYB3eCiUox2V8Bq5fw9a6fMn4IzEE7YZJ79gsdFlV1NStc86o2XUF
MnvwgyQpVVjreY9X3pprfvp6NI9vsmPgVkQiQxbyEdy52Z5zAaaHkDYjH16QJeU60c86KsEe2YLK
Am4uHA/Lsj4g7lu5BhMsOjQJYsvHPvdxiCFUzPpLgze5sTiGqHDo2HZoKeqZ7GMub4C3OEo3dWH0
Sn1MzoAO1qR4tyxF7wLQ6Wh82A87cqYRiahN+/f8159uHz8lBS36Exbc4uhfwJXS1/Qqfwj1AjXv
5a7mzqnKT30MdLWxJszdOrkEAlFp1wEzmb2kDWNARKIfoccmI7uyG4Q68jXP1I2d+Tdf3jh767B+
C7hXSIyWRCORbFdWlpL79yBWXEfvCIhPA4DAVhryLQk3EQ5UOK/11FACc70GQM3rOdj0PEin1mc7
x4rCISAAlpa15TUOLDXu8PquAcLvEYs4FD4wgQSaZTCpF4SnA1y4cgf1HixJof72c+iQESfDlCy4
BazbJ+sxZVRRaC41lnWgD9/hnM8Bq8dnxZS/kGAV3LXQFOgwFuFFFwXyvrlH+aCRE5/bs6MZmdUm
CwIuO0R4T6pHF+bgLGPHVmyQbqyjRVKJsC0QavtBvROHyZUG3eqnF+PnUgB3Y4fXivBc5nduXaeR
K5zszrmzOQ6v4Xsp0ibA5jVza6XzduLta4UsKPmkLGJjxQOh+xo+7ClzcN9Kow43RSH0GxmHmT/8
zV5P6rM+ZH5l6hWgdyfAxj1Qa/gWhBh6lFaH/lDyqjhfyUXlDskS4lWclKx9CthRjs6YPRLg7aAn
6MClpADKbPVibooR2ndkKSOlcWmMLbYBMrwe0TeTEn87fNdG9Q+gaJPXgCufAGch9ja+kXZM9smP
UdhpkF5p8RfvV53ibfIZROvfF1CRx3khdbkhbaJKplO4Y8GXdIXwUVbc4ho63c5s6ncwmK71BX9T
Sq83x0iGyKTSiDnXMSa7XZr+G+MEUf1lF+lsSMPcQN9Y+oMtWQBdzvuaEkxnZcH9IR7+4Zh2ZrvK
i3ovpNO6KGLKzCHSqtRpvlV/bsmKx0dIpSmhumyazTeAAfqDfxTaCbd7zQIEYoO3zPD1ZW3nzf3E
Fb+roWOuRiCzbUT/L4xNn6p22C9K/5KaqGRqL8THMvMJ3qcMNzjUjB8dLdatxY3CYHAUde5LDN4h
/BDi73LoiWsvjQCScAcQrjqKJxq0xgQq/jQAq9/OnRGMgUrVRkpciOgVjYF+iGTLj3r0X0PjlDkN
MZObjmRL1XENJYhfFE3bf3UXCwVxR41MyCazq1n+kmQKJH+1qKXEa7jfABFrAxdAkKlxlvbAZC/1
HFlsvMTSqc/8OKu7DskPb0VjPe9O1uqUR7XpMhMoLhlSPoP+UoNCWWzVi8LcWIpwvmqR8V5avroA
JoiqihWWEONuKLtyf1GGyX8lWyL+GxImpCBSCbBk9Nc9yCRrIw03z8L3F9DFimap8AaB++wvChLw
K5F0Xlwm9FbnC9HqkHUZj8H9jzV+kzOg5cAFZ3LCyt13Gco7VaCurVVav2dg6gg/V8XbXUC605Pb
GBaBrx1mki9ICPUS3GshlG8nLNJ9mjgahW1OKaXvn03stKjHLCKQbxST9aKT+/x/+2zIlzFCmWUx
gnoM9GBqyLasGRxVA4mJ5bGntn/ZsFKuqiKsVL7z2b1UG+4IlKyBkgbDnFdEs33GmAKkvGI1t2TL
YcQY3ReRH+2iPGXjOXX/nr0JgjbMBZwDvWn+40LkuCKWssYYmcBpMMppqyMQMJWxTvaFHuseHWyM
9uX8fJQIZ7fCa88f6quaUveL4xEtVvm5N6lxnpaIcgHH70SZrNftCHBHhPcVHScYfvZb7EkZc1lX
xqY6r7zT3MOkb+vsF0W5WpI02N9QuYHiCK90WfUu01LbnBNPc4wwPakEbwdhX0ogKg7dLQLNCpdw
7NmjWSypsvecpeM5U+fi2GX8K1M9qS9MjPgF70yO9ZZyJrhdEW5lFuQXUw7KQXLxUtm5j/qIm5Fb
yIxTLD08lVjirA3uDXacyf0tZQrebMZMSzMO2MVjy8zOdpd7GkohndcS4IBpiL250nycystrXSok
blxzogAmFeLpCPgZKjcDFPfRXDfpOGeuxrgQjM08LdzMaRzS5TXzk5gM7HCxo8Q1YtzQ8Uaubg1I
dQQjKw7WjFKk6zVhVqnfo4nIdVIfQdQO7RTW5LKGrcB2iAiZKXrzqMRdjuPtrxmZv+tl/Ji/mjeF
XYFFJBtyBdsOxceU3qio81vlfOdzU9/EWeSd11KFkPmDQpShBWYSrfHKqujrJHsA+i7BB4QD1tfN
wPBduSeWp8lfJa/eGPXXEmysb+r/Yqe5drpPk+W4Qfmp4NQJpyB3IeD+oDjKOQaLyp+mEa2Gek8m
MqV2+GZ0BAjPX1fxcSM61S0SVlv8ZXwU+CQ0Gci7JHQSBIhuosuzwQXFHFOlG+xA/m46d/ubVuv8
rwPKclak+ukBcMDl0Df3Y9sU3qgEaTcVTO9WFgbXNLLvug9KpvpMIjQMI7NnbrtFsCPjS7hyBW3H
qyyCcrXKxE96XsD8hifTES6GS5DXSu+Qauk8/F6OeRVFRz4wIXMR6iMxQoKAjBMWC+hArpnr7DNS
aymVJOnDociUzUWYXmivz37nwsdjMOFqyqSoWmFEY0PrM4iM0e73pvfOXAZmRFeE96ezyNjiq60y
3EOxMt8qzxewNEGK1v/WSVNv71+vIQCHm3dGz9+/j/Xc6aHfcBr8NLT++fKbiQwCIO/U2WImv/H0
FylgE3zD9v0khvjpdLuceva7MS7jhmqbP5lV+oii5C3u00QbgRFDAtRcS+aRj6jG9WO2dIfCMqPb
SXI6vqKHeYrQYmQZRdB90Y93riqEmcVtiub0Wgsa1jc0usjE/H4T2Y1H1Fl75oHuH0n9P7gZeqpr
e432aZnVmNIVbwZGqhvEZk/kTClKMx+KkhiuyUYdf3pw/HPAoSQxPIvA+TR2eTtJWXjgU7BCafH0
q8PTq5QtSNqT+1lFvq7bjwx9VMnPilp0DyH4FpZWgSpsw6ls2pTITK53nLpLXluxW/gx3Gevet4d
hpeB/Foa+Haju4OzlXy9AFSARaxlK1VB0e69aLHa4sE4bzV/OixFXJoirNEj52F4sh47T9SskVFz
+HHhwH68puSsSlu+THYkIMrg1lRkqAgh7fq7sWkJ1kXWkylgoBGkxbVqgnbhe7aJKGVuCS/j+BzT
1s+fB6YD632xbs2mMu2lCYn6sazcYU/bI2EEUawDrdjs8vd8Nx0fiA/tK11tqQDq0EKXwMxQs0yg
ukm6sNyXrWnS5Pc+EbwtuN3WuKf5Ht2zj5NhzIvuf5eIaYpq2dndlfCnc8I40a8dLr+6McxIJM1C
q+CfKmSHpbl15N1KyQilrwTW49YPNZyerv4tVMsgHh8tmwVsjzy+MOOCXvcutOpD2EAeJyDJFYpd
b8KSGkSjq9DlE4YOjXTOEVqjgWEZqWrQrhJqJRv/2LfiYpVQnvowrQ+H7/XQL992PEZawr//oTWS
0yJ69L/RQXoJJxV292azPPmi8+Y9PgLFALYUBE9UwlX1oEzhPzeb8kZs0Hu8PD7/Hxo3bAtN5qVS
KhrRcIuARxp4cwVB9NuVyue0WCYuzDhIX4nCR3/kCOpxdqwiHZY3EOX5IoZ7vKkqrFIJwxgAI+iW
SE7A/If2RRUtKTZIVlzfzIN4YUTcGcbxSyCfWiOl4kTZGpns4AG/+8LypaNprlO7uFKGCM9BLCx8
aNYyqeDeacXII7ONmy8fqvWpueRl7keYNEUsWoanxOws5YxUFzJR/YCu7xevO8ItYzat5K5Q/CXQ
Zbz2JPRMn385IhbFy6lW46fhQBWCqjt/+4K1rkGyv643/HJohA11vXtxZZYIiKTPFWqzBpEWzzJ1
UneocwRuC67ngCqJv3WLPEf/oRu9B1GXG+lPg1cnbeDjJoxyjxrUzvB9fRTzX/5urVRVrNp6DbL4
3FhiqxOmtoOTb7KYArEHM0nfYzZpNLlp+tlRDhkM25g4jpfrvebyoV0nXoP8w3Sz7J3El4aX8ys6
Y0sWLoXxPuYrA1rZ8QydeVvJVdwKcbajhLcn/TNHCetO3vbVMPH8evqZcyKe1bn6q94Gk2vzQtV1
C/EBVtObY7mFCGH17LYpbrMpazVFQI7Qyg8MIcUkid5ChUh8WPMhmqN0I3436w3RX7F+lU7uk6bW
TPAVY3z/yWn0OaApFbx7MeizQxqJrY/0T2CYVX00Dg3gMeITNaLuJfPZdUe8g9qm34r9KmEUivCI
K0W16+ki3maNo4UdBN3kW1d7zMhEgel1cBGQcrLE4xy7lXpj6/kj7OnyCsRAPw4thTurRPaAiDq+
oV4BHJYBkcfVKMSHigzman+vi9ozss2V2N9ZDR4+7C8+OzlrTN6/UMModGrzfGNOaHakLZchHFQm
XTgbKs+NgD0dpYUWbmb2lJDOOoviTgsf+08zSBzREpETw0q638gEsaZxQpN1LSdDAErmnQ9n3R6Z
2sfkRrboPmo0J/9Eliu6rfheKYeYKvtHS1ndcV9J0nD/1odOWlTTeB2Qju56ButlVrdzAJmPGHo9
dHQ0Bbb2X4t3jxs7esTSonulflLBgrIsuVT6d7N1eLXUPtI15ixZu4klK/HLgjSnIJRWqzo8y/UC
GkujyfcX86WjjKyKkHT82fUMl3qir7cWLO0ylTxbct3srOrSIWuUprfRGoKbKQwyf0nYdNUd7lAE
1Rgtz47OMGUpyDgJD9jV/BNGgPiW3Lnqr+D5b2EPzmUavYi/W+7FfGmPi90OLha1jxS27t0XKDA1
gWb8Zj2fC6soI67bmMUZZpQG+/eWJSuf1MyLUzphI6q5VTu1QlOQevxIFIqHzzSj+9vBHcLFS3xe
eIPdUB0WwEcp7fbf9jTBzahGtf8EYe8J522dzzkmqE4NwQIgyZ8R0OwVWiL5qwqh6a7uk2m9Id0l
eiK6oVzfXU+0YnS/noK5fJKjzlcZe8shjx+zHq+1yhoQD2cHyXudX0dEU97eIugxOoR0Ec2Bd1sF
g4OqrUqrdoZqh5rbINv4q6AyOLmmeu3om4FvxdJmPmo2Uppf/MrXPmUgdPlfKyjL6N6NgGkEcgOx
h+2HHHBg4e7a+ycUZuwyy7ySbAeApQF3QgGCFwvvL3zasQKZN/qEkBjGibo02qpj11KZ9C787Z3+
F8LfXvlnpvkAl0N4ChOmm2AJHtoDXyG15VL3xcMfr+Y90VdHrQaxGpMsUPTTzIJYayqWrAWb7RWt
rgzH4sffx8+S4+hIvfO2vgisi9/b6MSxzPpPAm6lSFjsUHSwgFtYAHI8B21fX3pwa4ts8QsLIbmm
ndu5autRyxkdC6D/3QSkarkbFxatsJJp+8ImF8ovTyyG0Vn2qez59RKfJI1itOPvDKUPv6c/MWhh
qmmb3DFwSVqbLovdGlaQfNkkIfNcTnirxFTJrClKcn9v7F6xTHsGjFrt/8iBrHyZmn6uK+aLpevR
c+w2feaA0N092MloFjD5Pt3HFD61a5QXd4m5j/J2CD1dm7YwIwqtIN1TpLTDRSG6VYt9Cyi4JQeD
eGXXTriqJE2Q5LJyqVozNq1rjjqU8L57YYEdaWb1tCDd2n7o7XfC/SMPGSb8o32BqjsabrneDJUV
wWPTjMNj0HGIIGYX/FNpfsO0f0jAaMNkDXaHfHSCJGM//Md0XFruLIoD5h0sCzOz59mK3hEkuD4b
TrqlrjkXTEBUKto0uDVfApj4aWgnescDg1sDaNlTv9MaMuUB5FNUwAMLybVnC3wNEyITkumamcBf
Ic1ngHhSeE+Dy5ScWOPJmjkpxYwAwuFQ4g97Aak6eb9jtJOTLcfW8PNNhH1+oD6CLRgsOVTmn6fS
clGo3iuS3ksIekYeeXeuyv7FbFHoEfSRRJMwldeB2FdhVcsXGgsTILDZcWMld7CsKuM4mIoVI2Dv
AA69o4J0KwKMirq52JPRDb7N4ttFidCCv0C8uQAd6IvI9gHu9wP3Gb10YP/MWgKiIah63hWiRaMt
rJLvhZyGzAzQFDtOVocArf4plljshUa9rQAN/HjXPclYtZMIYKDCrYFhzVmkx1eiui6hrYJa1INV
D4JlXIw3xy6RjqG4W73VAkghGHUnw6JVMjIBPW0D7gj/MqotRY2/qLfHqsQl78HNJbl0d9bZ8PIp
0kePNSWcM8P8CHsy9JcMiVWj+Lv5r+ieieL+rHexbqCfoAD5qIVab8/70rcUmXt8GZqCn26XCJT8
TVtbaGailtM+iwYKPD6AkR2ZJTmUwGZ5oVZkc9UfHW+D2zwOKXynhdGluTmkTEgtsihfdC4xMDUi
MrPNx8l/VihurC8sPaRplA+cBhfDEKoNXOfCG1bANV2OXI7Hv4rfAKBACBhE2knbTR/XPrSynCQL
CaG8bD9XeaQamnstJlC2jCuejjv/ZM+z/hB84hBneMGg9IegvJzN0VEVVmshjxO2aeqsjZC9iIEa
A12olHD9AVjSz1IsdqlE+nr/pP8V9bn5eY043gVxFDs7ag9noK4qu/EzmsqUHlZekdVnDHqgRbZC
ttRXvwGS6Jj4vUdaDUKheQGBww+W+r66PHzmgXbWsgFtA31KR6HU/iFyWzY4rXnjh917uD381gZJ
iCt8Svo1Gwro16AJfKWwudnq22uEEpACgHjPmBcLNuznYxp/wvY/Xa4nIq8hUf1EiDttFgzujNib
wk2X+0Rw5AgPDrB+xkYX74pLvgcrge93ING8WFRZrVXQhTYaq9gjSzxQt34va3+/rmG7qSCXV6or
+5133pEGi31ZrajiU81AEVtBpIHESUqrvUxFDZybRwLgFqKbzMbHgOG6HFTtmjYFPkfx20aObMbY
w4CDTBgJYPpVfOgiBAr/Yq+iO6hxjqDINqEnjpU3pzGmfEjN/Fw5Ny2KoncLCKEZ0qC14zWr4Dho
3ULcD1nJXocbe7AUPclxQmYxPCqfbr7lTGamApv0tiOGayWmToS6EBFVGSXEtYqCNeV/x9kUMP/B
ipfM40LUfcE0lfyff7Fw+KMaYzfgSO7Ne/Hspeygf6oEsngJeC8LPDBZOMJ4BOiQFADVYJLa93xK
8GBjmhDdXzwbpQ02dOBFMJmxJAdY9fWsFa2/WQbkDnEXUE/vUVeUS9Z8GuW54RpjNssim/jkrvzw
xOaqiaHe/41VkENy5Od7z+liPL4R9c6fB5V2TqlkfRga7rWcRfXjhsXIAFhqLqx6fhkadZ8ax0Be
oSxRgMn8V8rOtLJ3e8xPMRMdtVQLanhOkjqxMHSkmCIfAECjLTGjVHEt/bpvlaZ6KOJlYDAMIu+p
O7HswzJtKw0hXf+OuIgy4pXii2ft6CIj3tzgMyhVu8klU9X+dXUaMcNGCgbYf0/eaGQWGKt+bm+L
qsyBflDyczp+2vq8MJAvJd370+d3GjUb8FQmF7yZ8x3mbt6wnW9BwZ9i+FzE1MEa7baOGqmTjspA
ovSPpsfiLZFR1y21Ev6hXOmNXQ0LS5bdw4CbZwAkFZEC6L8C4Mb1QO1Xb18ZsOPVKZrqGyCbC15S
jTrqMU6wKN2Nl1xc5LFHjLeUgi72c70AzgP2/hB49X8mjUsOI3LsiSY/HXXPBLEPGZKvX3yZ4GW5
fyvwfJbMeDbXD4cPlVy9R2bwMP4xFHXxraVHXSwIl91HfupmlXxrUTGUbU6GJ4E1DK3qfvuK/3Cy
w2YfXJwHuluMDp7WPRodtRkhZ3m1PixnbHBhSdzAeimtTeX2ex1ZwnqxWzDbAcgcJxqIGKLpPVQ3
8nMbD/rrD1fBYR+FO+E+24PDPAhsc2SJAfIjTitY7yQVo2sBjEkKm/FsUM87kEshBAES13t/DozH
PWOB7pJZ1qlMPo2J9edvv7gALhja9UeL2qDrxi1bxeDzfjM1+mqgnj6kVY+jV78OtzsJANlHmvUf
7bNWjAEmv/UXRd7ifryjikRoF2OYYbESYjegvXLmw//d4V+P+KNda+Iv+p1HYeQsfI03yTZGKxCt
QMHr7XVXAQ/DCuG0L5ZJ6ScmQQEMGxbA1BlECyjt+pBr10XeFe8MMsF77MGlvljrul4cZpVvmHsd
A2kUkMsNhzj+K/jnsVt7NEQ/Ahh3DHw0HcEzQZ3on1X5l/BINAJpWcNanFmMOeIWVAXrhfcEZIE4
GbQwNLSZ6FqeoPIOdC93umlwX9pQEUa4CNgd/C9NWDNRrmtehUO72xEyre6Pn2rp/VKTOWHEeT0O
KcVx1Rk1lnnqTjsKJRP+J0HhgZGx6mCsfjnZvUEMt3+HUScIdOjK43UpsW+RtCF3LSkPxhCHE8VB
Ti1ltTghb+R1GhKm5dS5kk8iLSsEXAtZySmhO1kaHxO9Xe9NcthwylGB2VWxb3xW0i2QNdgOQtIv
vduFg8GTG4uy+IX18acxWHpzkCE6hJh2AzVfngo50HY8qmgcSWQ+4SeSn4zI94TffsbDwZYBBaUT
oqcxmdtwQGKJUsl7YoUvSN8nO3ooHr9HJvEDK1uLwlig5TI0g6NCNqh4sPGdUJFxM9LmGtOnIEDW
WjymNcyMtqaq35URepFjSRvgmT9s6sFj5r81QueXFkqDuigh6PXvZEGg0LZUjFCNXPytKwU+lKp4
wTOmYOX7TJAYsTdgWhthoDqUtTra/zPG/CH1S9MeJAuIkMTK1devD6DPnekOApBIblsy2DYT6qY8
rpKQVZlRsQrKWhu91zpdqdizxlaqJCR/Nm4lx385uZ9UlIBM6j0oIF8Ze/eHSFFqSSRIUfRJQ2Nz
ONIcLvnKn471KtlUvmTHkWMQ4xARZnb6BSHe0L0jm5Qhj4aytT/5wn/sgs+gm9kAATQf3e2+RiC/
JvTnNgX3HhQGsJUJmhMFdAiXeM77LOy9UkI/B4ffKboeNcwnidmbznMmP4RwXpMw3wxbLQxGSQU6
K3ZZwBrOkbH/t3Sdo0QsIlrMmJzu8t26AJie45VioFSEmMJUrZH8gcbIuFaDX7w5wAkSL6AlblUy
sNrIEHYin1HYavDuic0Ghp7urFzvmUeAhwiHK6myXY1tFt5Pzj2dnQglelkdc6Bc2li0rEfVuBSU
wTZcnwi/XD6s5+ao4iHLwBjn2kyvUphKbGjNmZ44y50c1yK1Zo5xJrLuVKjF1L1SEPlXI58nTbS2
2vhirn3JbKaikKBHfhlNEgws4zYSK4e3OZTrCyaBtQQMRIwy49Jr+TjRnd/3FeFCkZa52aZb7i1l
AnPshaUCEtzad1H+uC2NG3K+FM5v2Jwv8d/udhc7Z2zxIkDohp161fnqAit9gr5qBNITlRLi9hy9
MJCGE2Fj1sdXQUE4DC60pP+4wg2Nc0shavdbcfFvLThpG5NS4jMJaV+hR03JwklzGiwPk03czt1i
gq6nvkLc0BndzpSGnUzUiGkH23rSH5jy5ocFRXAu0igpN8hjfXDEmBxS2PYU4vkgj4LD8hNZnO0v
yb8kis5NHAFBiILEWdIkXaUdSWL59QKvRf5ujGGuNwYIxFvo1CE5+LNYgbramV4KwNMMMle9Y6hk
0yNPQnDUCgsYIKP4KI1bGPfK1qwWHav0LAZ6X40b1j2BTCJhnro4U6P5a/ZZQzaMA1yT6s4Q9xXd
NHf9Ok0Q6wjk6fbhp5yfU9DngGNwFMNHS81ucX95328Q0gG5kXVRMhg1UeFyGiPFq5GlQXyoNXs4
Bal7alvRNl4t6ZhJm+mWAngPizvjfyBhZvczSO406rVZ/LeW8PgvjP2SZaAFdCnbqfIhnhc2oNRi
OezjbyT6tnrUJ5ho9yqewfu3C5Ha92QTLSk7CZ/dIWprju/3ovPULmNimlCd7sC+lVNA0D45SFSD
+PTpOlaiLIifwLVXMUhQkeHIFviuAYsPyT65R9RJbB/ZZW5SnmaQ999fhCeRt1d7ttjDFcyrG/Zg
CbZB7PnJexZyFAKCsHxVfoo/GkJfRGLS/pQ26gUzUu2qpz5I7KD74HwS1mCEeKRd7euMU7A6sWLe
JqbWp/Mu9WdNFEMmVLRExwOFKP7VJvLN06Apl1D4VPEI+goaAyYUQJkJQKvtZSjzXLtY6Zqzur0m
VlkqXKBUBJ1sxoCvxy1ESWag5UeCOYoxhfvZ0IYMd/41GY/iAp1vCdL0cixShtFJCoiirOlBng4D
niGwOfJDGnTH9nXLJuTGXoaMR1BXZ/T/XBnYZ1LFeoxiUJlCizpCy38pXa8ONJfe9zKhBxFiTYH7
LCvfINeNfJBrneNGSFXvW4tVKgd05YK0px38Wvaai/W+NNPklTTewljYAjUx6+PDy484spirmjRK
8oAX+PpzHqb3NS2oKJCpAdPGQcjdu1q94E2Hn5NhAg5gH4om7xvM+yyU2GHGRRHt+Zpnf5fpdZCq
m5Rx3v920LIftnQoTWAUbT/O2rXHfg7PbRtx/AYWiQoUA/DPx/8fFuXt+WrCgX5c8gejEFq5rWQc
IlkElA4DxvOSvIhLhI7mRzMYm57DMnhplTOlJ/DZHgbeBYTEK0IIWIg8Q7/rFfKKXNLgL5Xwd+tD
2mdpWvX44lML5O9DtexYyLh5Ow8U5PppTluOY95FpY/XomTJNc3T7ozUkIMLYi6JxtyVzLyPoGCn
eo7NeyvgTutK0cm4A2BAM9QRDBbgdUBHeRF1cAsXeor8V9M3ujY2H8tr9yRfrUt7fFh3KR+F1FeW
eSfYI8+xB1VRg2k9voXFftF+AzBU/bOe5JAqMrveRvWOZlhEDDiFuuNXxRN94jEALfj5FpgLt3cF
IXRm0Ri71GX4Zfkx15OUnJm/ocNjOfqrnuaR9l9cu+clxsP8RHlOGTn5tJ9J/OkyPJZWFEDcQpAt
p4bCPt/NRts0Z6TwUB+LcwMkgVKGE4lrABl2OKTROttQJk3ycNvUVYu4L0hVgYSdc2BlxpLu9mrU
2NJLEWbaGbIWCdcxGpdnDZVl9wJeDjk82QeJN3hnjqYdK+MpLV2I1vpAC9ZAn6tGSXA0KZEE1KMd
+vYaAHNusrI7ooZGtyQpklvx9dBo3cUY+qjGMCZ0n1EZd+UlTuVJFSjZOz9KvGcMmvdnrJisRalS
Aoaxr/b/Vx8B63DFLX9UESepCaxcEbLnjKKTbQXpC17//97oY2JS+sMmSUJEZ+Yvz9CXnKp5k5lB
S/y6EyiWhtvNsCHHn5ATZ72MFR1ee/HqRETEBzkTzBA7cCpfuhAGNizHkJ7SApSlny0F2kBFjjaJ
hniST128kseh51MF2JhC/WVY6zT47RlvK+bnJhdJGGo6NP7EEtmtgS6in9+LQCwEVA1RrP6lcKSJ
tOxMfDKhFjV/W8IhFXtnmnRyLC8xBMQfE+JxgUrT5vSAAFei3FM6eZSIZGBT9o+bjW3n66zI2LHE
beVWCkRWe0IeTuiqZjSJqT+YkIr4BdCZDU2EG7hwo5wQsCsSckgMR0hUD4dmWkQ/BOZH2Q0Q12VF
cDiUqKx/SOBPpdsDamykwuY+Iv1qDX7oVEIAUCTDBqQMi+KxK88Ls0Q0N/6jsLmVpc2lLMiE+tGo
CQM8e9y12pXQcP7swD1m/yLw/9IivwknSMwP4Y6Z2J3vrPx+G4VpS6Rim+7dxQrBTDIUr6pGJ+rI
4xgNL/zQm8LWAmqC6Ixpkh7RHQda7x95AByQJQoIxBO49PyEL+QTVLrhoSQalB+dWmdKTa1ZmhbT
lss5WN5PEpwife0NHKbX0FCV5fJVOwHXm7uW77i7lGMtkAk0xJbk3wJEm33z79bOdGgT+gyEOZhF
1fBlWY8l0Qm2K8kurRnYL5MGjI4HpqNlot/KYBdFnrzxoJAwLIxuVkpSOYGKlS1Q7WMYIJ5ZuwAc
Sso0QCF9AQpgfeutBkJgLzP4qT0hoeBE5XwnNfTE7/2a9B+MXWvivYk/n+FWcoNOwuimVYw3NnFq
yzo58LC5Se/P9CY3E03oKnNjjbnG4SQCRK+d7p2ur5Z1POUmb3qzgUFvvULh43jxjOU7nEkiOiGc
AiBzjHfmQhPoQnuSPSWx5IiPpQvbC4v5DMYH0+shXbRnpZ4HE74DZMK55PeJ5toQuXRIkdpyWxNx
Dbwo10jQrHf7ZqDKrWlz0wCXlqNwzpXXkb1D3y6Ce52+pqAOPtTjSe/spwEOqlDxiXKUZmYXcGaM
IvcBx0P6+amkrhnD0KI+vXgwLbvTpKE/eqPYj0/vOl5DR2xnQztpBunJva9kPf87iurAX6NYtKsI
Py4K4kRViOZZV2sxbiwG5mrgytIOwZlOx109Px33U6peIjW2fYiZ8o94rxM4N1fzJJNLsvy/3UZO
vrZ4IFQ4qNa4KZbO02PxXYpT7sepzy5hoEIe+oHwqCIkPbT+lxebMJm74GhkUHfbxMv70LiwxeqG
UFOUcUmSvyuvcPj820g/2SNjSFPMdEkyFUPluj8FtHWCLpNMLhxMpvuGYsW1z1WQTpXbfiLPUSEg
N9poR9y+UErimUVwLJadc3mY8aSXS03YXJ9WeaEY8a7IFurTfjzEYDH5dlt7FIDAEekE69cd65Xz
+PmqeiTw7JN/t/9tvCnwl41nbRDG7nYvkLCX4FkDbiUx0N/2R2Ha52YaWFSpDN3EBOlcphrASj+9
47DOud0bii0bC9mqiRefBtdm1OA+Zyo9OEQ8wsXoaFEBdfqqP2kMT/IypFyI7SdtItKkcJGSYeme
hD5LW2nGpHhnDFAfIntYBNvV8sNVxIp5ZI5QTQSHHj+Fn+6pgaB/GnQL+YP9jD9k1qVnmfSefMFb
rgk2c3D8XpXxk4TFHN1/yTS0MDGZhnBxqglz09rLWIdhuDxlTVtVQroBcfLHavYlLrCExg2PxOPF
WrwPtK+QSpCsuPb3yk6ahksJ9rBoicqejJIQgJFsos8ErO9XKIhPQIeutpiCaWluHl5uKsFFfbfv
RXg+AHaSdJ/yzaC+6cqjNIr7Q96rL/MwDck0LtbAAsqzgW02P171XhFgVDpCMhTCavXIlGbQwdyD
IZCtDSxQ02whGb6+K7pbG5d+hA29t9r+LwszQtNf2N+rkCVrQ+LyI/vVicnJh414MOLW4yND9Dr3
bZ5s4YFy7DF9RQW0UtOxrjq4kzDEAJMPWb0Xq0Oprbzcq9WLQPvBSLFR3l+c6UsVCjhZ2bEIaxG9
33mEjipAJJIL8+Qp81fiqEQpTYSvHSm8axSqz6V+QSnj6GZTom29xB/ABZ7dITSpII3dRDl09EnD
120Mxcr477MgSzHnLZaSmgRnfp2aVnMSwdcj283fpzhUCXeUC0yYxPyzHeKel+RyTBnZ11OEG0Gh
lPXpPjFncM6Hy05Q6N8Jp49hbuzMCcMYZUp5mvaj0jLhJ4igzjlw1uvape3LPjRCe0oWOCwX8e+N
5EdzsHkQ0FL8HGZg2vR87fStVvVoNpptt1oGqn6iF1e6NkbGXJDggm3KASA7VVXSXUuepakCBmvl
6bj3BFsz6iZEV9ev2oDP1IHMBQY5nu07X/lXTrwqryXpJlpqiiRaSaGExZqOeyTtiVGgMzvUhL4l
c4nT3KP0Af4HM9QWyJgqglbj+9DVU0LFtN4MQVzx0HqC7AXBtGWmc8eBWpAs9/NOxZIugSyo7J4N
QzcgurNtr5Q18+tECjad7jj/kYBZIBEJDLd8QNS/T/s0GZpV0dd5vxeqyrXX+ljnDppicBGj23sS
K2pVYmDMpq5Hm7aGx6zz7Jsf40kAgHtkqj7Kx7OXj8YL7qhEUn8nvgaq+gfsV5w84OtY4F1YR6PT
lLsCytFaA7+HP81Wg3GHd2KezF1e1fzd7GcDHQA78MLuC4gbleUtFBFnZ3dLzcaxjhCmCz5SLC+G
qVWJ3UauBpwiazUbAdJqY8e4ZqduWaSBFSv2L5MjtVEpNN0OZFnzRwXnbulCu8L72Bx1Kri0lV1n
ET7DQnWpmQKcQkBEvy7MVis1aZNLih9R+ahyK4QqlRNG2FtwqxEgmIVsVvuvYXaF6CD1iwwcPNAM
yit31mf7gmYTIH3aFtIfR0PkifLtiUFNjN+H7dTIRCrEfcIH8VbRiqLlbaNS3XnGTUL7+fMSJxMW
oNCbuBauBJy/talwmIZYnwbDbEq+xnRMGrj/S5gTnvCyu1d5yH2pMzZUpbjN8+7TGDj/kk+Lkd8W
lrCl52T8RnJvjKbltBhFv9JvGHps4I2KiRocjaE6zzgLuEcmocVQPGJCCQAavHQrtcKaEMGM0AU4
/V3GaJbWwtIxHqDDnZki8Gc6R4FShmzFtAXB8HDoXgPO5WJP8V+w8lFr2VsNjaL0S8dFm9MGvnAL
ZyIaTV4bSBsb2Y2mbHW8hsTbo6D8lUhdvEWCQQlZVi7WY7EjpWBjHTW+b0x9a5E1lbXiC7dG/m+d
GmCbEsTLc/GZarxO5f/Mv3qulMHkF4FvyasmDsSeFPQra2x7OiLckexS689FmuficOJzyO5MQwSX
es7f7OKluYNi5y6PPaQ2+prIi/TeCOc/74K0VejXFvLtOPIbXbD4pz1bpQl6cng+Cwq+nr3waQs8
jH27m5yQbaTbHX2/ggBV3PW+z5lXUmCfNZE7SWJsCEX0wmtuUkD9qg64BsXm9shN7+PSDm5XuJTg
NKQMAGlJQ82fo9ay1W0KSMSnvso/dK9RLtz7jbq7pEQFZVtgMe/3auVHjInDkDmx7hbUSW3mWCAY
I2rK2NTVgzcEzGzMYUh2/rj/OL+9MAap1NyhzkEbSfP9f3RXvMN3pLwTe0wcxiIvV3v+vedP6Nwp
8z0XImPgJYqR3S/ImfFezU+FqZ2xBp/7UqLn4NDUV7IT7zJybVC0t1Zh9lRjbvg1jaNRwU+/AiVm
hPvmx3aCxt3HJtzlS9UhFAfyYKjP7uBc9VDZ/Is0dyxKCGkaKLiPvd8T+YjUGpRglS00fIxJ4GTx
hG1AIo02C8aNSQm4WBkrBXb8Ie8p5m/z3TdpjWim5SMuJaStLDRI8X3ge0m2WHeijEbqKNNIUoih
mCd2LxZMKKDl952cZHZVwrn8d9KHsvLQ3Le4PLYHrVzObr/uq/JxRrc0l7HMYnGjE6QUoLG8lceP
wSXZS4yQagp19lUp8M0vKfaBOF665NhKdKQDxHOM5S+YhnqpHngIY2qv5/r1Tt/ZbwcIaBaGvO2m
SGlqORcWwqtGwCiA8QMjTN+Kd63JHOSONJZA0sJMf/jCqUkh79absglPmbAVxn39cSy1soS+rP4U
AMGMen5oNgBrFu2q4LIMK4RrDFkOD4lUemCEqnemeRsstu9N7MReRu4DQ+Kj5zLrDTj+nDTmNxwr
IX/8tqA94Fts9bwhn83tOKYMbbscLBYkYhbJVVt2kp7SRJSm361Xqqw3/0/fzN71vKEq2K0QvKCv
9LIJtLFx+VL3UrqnlPoN5eOlBjtUUJSwPTrWV8eAvdHHQDr9ZRGGdapGSI3fBKcnWFV74nyFMciN
eaoXuqHprb1cowcmMKrbrXM5ZkmHLBaaHVOfMoNrFAOoqg99um/W47w3ZGz72u2O6Q8yMywhP/CY
KoXPiGXsTQrA2DYhFnnZrsSl+T3a/4JqALw+GL7z9OE6NcjBez2x1GYMUMvD2WaV+UckyR0YPJmg
6sOc2/hvEaMQW7x4aWsOsqjCcW/mlToQYJk0Ndk/gkTW2/EKRzbxEU3QqQVF4ZfN1oUEvBM3wgpF
FIgQJqVXzjjSwbgvW9eIANOnof5c5xW6RhHpWNeGtS6ip4/dpt8Cn5ZtrRR9Cn64zysuLgwZVDiE
nmsZNv4WrWOHmWQ1s3dutObEqOQAL9mwHcP37VRuDKo5QeNMO/d9G/alkWk7geMMoACO8A++hr3+
F/EvmynysEaPaXFRdY0XymcdwjMeqy+TnkP/PS1+Zw+5me2tLeg8NybNKYKNjnSzl3z8fbIB6q2H
sSwaSEGJ7q4PbJ6lncKvobA7172KK6dI+V6x+tkdqluO8AnWHfHSHtUAxnK07HVpdIGJPhaxmb+i
sEHbj7K7byqpgxsuF4fwT9/uRPoSB6GQsSLUmZTnY7jmpeEFah6sKbQSGteAAUfTpZpldYyVhIna
au5Y74p3pnKjxsRHjc4RBLwyllVBOf4dHuyBFdlosThETmEN6wVSBT/mkaMHzxbzMPS43Pbcn4pZ
3bYhWy/hRLJ0wgdy7YuPPxGU3DoxYTe8wprPK8S/aNGBdnukuSJFzyubAwyEzr0bjTsTVQDff63f
AQgdmsVTWqExqMAssKLmVX7R1qG13tGp3P4DNdwXCyVvJfNbazI3gWSXKvTpqsgeFKYhgogAbWym
DXSJIiSAslG+LKkWoHwGKWt7pSqceU5NBtgllXgnpY0FYCl2RMmSsoGVPA1LY8hw2fgvPR1enWwa
fyl3mDdxBTECqR8ssDdP0lXmREKwIy4anzhSqY4UZeuuwYV2HXKgGxF8xRkxMRvGMS3bd/FLOlA6
EkIq3p+GwznRe9kMcHnAKVTcDVcGW+7Ql0L/4PyTX1bo+vPgFVLq5VI8dZth3TexVZEdR6PEGaNj
0jzUEFEFwSyN3fr5NGeBN+voyqGMCBldpLANbd0+gs5Yp5qSESHbHMlRW3Y3515H/SdTvp5DrxyC
9xvywQnbXLUoHcUm+KaUGNDzadUYRM6ZzhUf4A4dD2j0rLaSLn3Vat8jk7i2+BDN/RNLSNqBkbx9
rkC/kjjD6AV2FUooI0I42InIsio3bIKx7dOhhq+C7GOUTCZODqiY0/zXGupSYRP+dicdoR/gGMPV
GNfGnBSiA1Pr3yCb6PoJvdsvpqfxpA8O8l3Ujh15crhx62tkWh+Vi6x79q9K1jrf1cvrRrOWO2UR
3j9FUZsvMuDEWezWP83VaxsWuUOrBUfx23op9aSM4jCrrkkQYhrUeLnAFbYEtr3qKXaWNkC8e//j
piEZvIWV24KNZKZ8qybbEBu+0LKmuQWFs+LdiW9wXTP1iGJLmb4WweNYjmL1una0UvFp7SrRGDx4
WOyw7sgFJU263tvVkc+SBE7mcQro/M0es/DyIHrp/8eEdNfXVVMi8PstrQzXSSgQa0t2UWjNQVge
AMm63LCKlv22LPZ2a24HoDBY2Z6OAR0qrFIu44YVpAu7MDqwrRnEWrB0PdwoFqjXHfBnN7ZiQwic
gDR7P3gu0kq6f+Vn1QHkHZQKGjFAIQO0DmJl2q5HpiQm9NlF8/O7ag8GClR8rQfW7dGkkowVGZ+r
caJxMOWdPVrGPddXyqtoIHY4w4dfAW8lLMq4cUaXCiKmPZnywpjeWqpSsyrmWHv89U+krLx0M5SX
VSVaxYoBmId001V3GN+ProMiJ/D5fx1WqeSlIqG54sETKXM2qoBw/Ifgi7+9NjrFCN17Xng9XCgW
kV9mT4/oyYW6ITP7ZfZUdnlGyT0gJGwPHqTiifirYKYDItjGa8L72zjB2G+XtO2DFRoUVReOheDp
BIaBcF5OljEKPTVvc01/FdW61+sf6ZjNCY1TPMV/Jac+5mQim3bzK5d1OKSTHmxDQGYmB7EpnZfq
TfgZEyc3gBMoEZ9DY8EYSHwPjQZ4qrNvvWa+9IfZJiOFR2MF8JH8A8V4ag9yf3bimBwh96JFw+9A
Tnys2QAv4A5b7sin3tYI8HlE1Ue4tNOYklzUOfNlpveD+0ooQZIWn+L91zKAXqRC1dnjNKucZvDR
+zEAZmYxVpRDOnV2FjCu9i4bsm1E1lkc0Hx7iOkNDOxVKXShkpBUgQFtpAB7W96xVQjoR4IoWyrC
BgEagDd9kaZf+ZzaGwSkkM4UeXFtDVcZ+qcfGJNEF6XG+1ILhI8v7aU5j9zYcVVPnE7zP/lCKnHh
DrItUJnSIYpty1DH0+PEfxRzwIheCg0ZpsPIn92/hhGMrPTUSEfrIkHzYjNZOu1f6gt8GqWJgfGP
P8My22oYRAFxkmIdNquzggka1e/0ZVIb+YiptySKZgnpA2RUKlPLlR2+H12BHjGQQA65zlKcS997
gOucnQkb5TWaZTKHu7mrW1Mpa/7dusbAJg3KeIQBHW9eJmrA73FZ+6KkPlH2EIKkujGNDZfBetDa
oYXhR53PCOB6PjPWvZ5qXwrlv8rTM2EOhAyOSNSLWAtxPGxqCKsqBOwFE8T4wIJ7iqnawm3AF0eK
/HJs6fKte2dKFUxxEsV1KltyDcQhLQGJ5FhBHHEHuFPMf01Q27eG2FbJ0oiQizb4aPpgSVJqTGT0
khgneIpFfjbW9AYWnomLJ3UKlgP+6At8aBXVCOmiCcCaC7ZdpSc/1Yy9bdFwOY6BFU/9Bt2lfNIV
YOUM/0Dh7H12CiDNBrWwnxINGD+oui9W21qAXkYA/4RZYyj4yoeM1JSi0jXbEkdGIJMsYoVh4SjA
lPX1Y/5X1qUjZv5lq/6YPwN2etMgVTvtNmkPZEQnsOnjMciH7dsX+4l7msafXm1E0YA1KOFV0GwQ
dvPBwNADe6pN2ArDaSh1F1DOLAVXudBhf9rKOnkfEd7rR0yb2fz3OqzUVwWTpQSnfXXUUE5pO3P1
zmPxuMrOY3DjR22ECzXSiREzlTCo6iB7mh8FeMvrDOvAHT0p3yNyQ5xbaVFOchxAJyZIZ/mvTrME
92UI6+BVTjX0smHbJhNSEVseN2Ek5IDmexE3y2SRVD0W/5g0YBqbmBJErCsmgp6YxHSonIOxiWog
1B8Ml4pZX0K4/SiNmorOd4dDm15936y4RVk6Fg9QEl0+2V4kr6Zp6a5E8kGgTVYo6P7ZBs5Hmyfg
lnuqUww2NPhTm3Y8iUhG1XYsciCJ1xPJJppR9nQ0CeG64YHbY4HToM+yLtQtkQQnDHMveNV/kBNZ
RGs8Wdth8oEGd5WeJvzq5KhzKijfsLa88SpqzMRsqq3TfIvo0I47oE+L5H6MscUQImfJfac1+6wH
6+2yEijZP1g0AHZCLp1tFapJp1ItkjxwHmkeZa4X1Ofh/sixBsVfDOMDljvlsqiz9OJgoSBoR5Om
vPQvnIIDUUXQbMgG+atTH2WGYGsABW/m2lgQr2F5zZo+LDdl3bENyxbFEyZCPVDt8hZAAkOQ3rtp
aeSAKElwsAVWVmZpqGY6yUPDsUKQuxKlHLPw/eL4WFangV+6/eMv4Leypa1ffEZDGUsGZSCeHG+8
JNdJVDyFVzLskO13YWQeGB9DKjO4m3Q4i7xWygBZnOfgkLDxmLTtIa5I5FCG+1AiInFKbjXzNtbn
TF2r1A5JsG5ZxBaeY2NB04KZUWR6oHzGswKN4jVwt/u02GujOTMvYtrXsDhm5X21IuQVg1hOETTk
Tfxr8MkYC2wV3Ood+f/K1qSAkUHusr36NpDtIdCB3i7Qpn2GdmCaCuMxDUt/OrvtB0qO3q0BEkFi
+exeVHjMyJFT7mQfk56QGGOqbpfvz6716i8lgOM8NGXRjWnIwhRY5O12PjCF9O8sThk7+Gev8ldH
LAryI9q5PtLP3Hdg7aTvSn9mxQMKkWAn4v65c6xaT5FMlLlhMqywx0/vaNZAck2XWGvgIXihNp8N
M+zXs8Sd8R/DLtFEeFUtx9KqV98DGtN69Mj67MzPzDMRpsLJIxrn8wQGnWxbDGl85/ctVjyM6lQ7
j4ZDhxOaoPlXvqJxwJld9gCRaV+9V7kTIDtRC20Agki0m7YhtcTRsXtPpSVkxaZn1zipeMY8C6pm
NpWe3mW/j5DdfsuyhcYelDy4je49P+KDSl/soX1WkbF8fLOzI/fxz91BJPYvbbGdgO/pPSRrIHKd
K0x++03luYLKxrY321Gie4+BqWtsQHgfUCC70ZMsVRPHkL+hXmc70Yebi9Tx1EzzZDwDYxH5xU/s
+xCJEL2qNX1m0x0U8vsDieDdKJuo/j2ZzKZWvRh947/s3Cxx6j335LhkKOK07GJErxu6a6gBimQ+
WO6abD7Ad2tBqKlWJbRadkFFFXSVI6Sr9Nc9jpB8bIyjrnaRjCX57wBXU9mcXW0zl7re4XVG8Wuw
ih93doimL2fHol4VoGQtx3rA54pjJP1wbr3LY2liK1T73Xm6r3FHtTWlaAALy6HXYOYALIgqQ3mR
9rMP6XwTHNMzStV7Ggz9wJlMh8qY9QtUqfj5KDdvISZPOw85fO1UoDKekep+r0n7J8EOd5Mwfj8e
y3i14+YTI4TPfSA/yOri0pNg4ElkVnuQSl67JiWJEwh589iAHUkANKKKKo241g7BBNLCSxOGYiQt
Zw1jcZUU7IXn4qS/zzoC+8sJiDnOQ+xaz/I0Htsw9/N+ZR1G0+A0tMhWXEemXcECny5I9vHFDdzg
mwK17lX+OuGXbWfvVTETMhr6bb5IT9NZnT8Nmx/45S0kIJVUhEFHCurvNQTfDsKFndxOentCDa5r
RqHT7hDok0a8OC6PyKinbbSbZUnqq2ut23M1mVBlsMQXUbmxJavcz8MPkrWuFQij4dFQ9wNIWGua
GpVCgeRWBeHVOIQECZbvP/p7QKIViWAe3PcYIJuG3MNR+13FgSZAMgZemhCrZiUM9kCh5/Z+qoih
B2+m0YIFFKzORQojB8Z/mMBOHltVrTKui7e8pSHRDXjt9TSFe0HHIIuv5794wCFAPSjVH2wC+3Oh
s5tg0F1/EGYnoRpunv2wDC1Rfwuthg85sW7czyeBygvrSrNxZKupKKCe9a61uiJHc32x+IMP3AvJ
IL/VUmubCv+fwMIHwmj2TmYSI6dm1CR3F3cCGA2RvymhFa1nUzOsHUzXGm3+xXBklP+T5BNwNvhB
1N6mdjEKT4Vq6+su1sCxIaTMidjcf68mo62Yfy4MI5+A7ItFSupYdx4ExllNSUlhLhYFF5hR2AGy
x6zlKCJs149fVgJeXiVccT5ZejcG/8hViOerzsQTDm7AAv9ywKvkNSACZjUvS/IvIBPBGnSI0FmP
eLoiVdPZfd5FXAAR3VRF6j5w3EZxc6IZv5FfXdekPAV1mr7v8gu1czKakSbSyvmS6vOMm3SxJCvO
/ux8K6LFlhpaie1cya8nuzoumRH7NQKBJMh3MXwAMDO39xf4kOjmFOpe3MOmFo5XTXZF+ftgTYZ1
XoOzRN4Dy7FO03wSb6BuI0dUivsoU91yGAwX+X28B1JHfyJQU+p50BH1h+xNzhC8MBwgq77Y7A0H
xtUBqNW55jWq3hW5w13tQVbSpLvexXdmPiA6PnZteR3Y7ksml0Qi4nBMCqb9NzNeYvazokUtxsm5
sbaNFD7ZDZLmIAH7/mP+33bd3C8w1UqrNN9Ju5mSsfAjYDs0C5h9sLn/KLP/OcNXikfB9C9KGsnm
ryAwpOkoX//QlkBze0pRZBYYRDvpK3VFlpaTkD2ceRH9NWOsjw8bCX61KOwp6g+wpcS0voUuMADu
tf+L6xm/jxDCvjDM0t46OHM65OOuZBGWHkq+LPKRYKu+yBygZIMr2eYc23piSrIghdL5mwWN3R0/
t4QboTCP9jh8eX31EvilBGV4PpW+417nsK7i2LzqdxnQrEm+92sRmnUP7lKmLLwXst2DZQq+TZl4
3/2LvU28Em3cgbOVBVBHygtOOU/4GIq54IdItTZw66pmgFi53F+MxUik4bNnr6rNTBA216r/YTa6
Uvk6136intF9v4Lpb11WSzG5socM8ZO+2Ro6fZQ3WZ8FQ3lTFS7jnSlqQVoWvWDrYt4PPN37Vb2k
LT+N4+AsRiWuV54JAN73l72bOJqib7IIj1krGcqbm2RXHQ86rpdkMVQv4T8fixzLhEEZToc61kbj
qcQRn6tdSerqJUx1ajqWL9sxFtkkgfobsuM72mNNuj0eN8iyElIYBfRZYUgRhJJIWnzm6iG8pP3p
nwXSmtSzHjtq2wlLABds8V4entpBM0Ten8MShxqKlBST0P2hmlXqoHCPB9TjZpMIkM2Dpw3uR5xF
fCrNksNPMKh9pKSvwOJodMOdsdCNtWrv24/PJdyOy3xhsFqrFWpf7bfqgowQwv0fByUAcZvJT4zR
yc4q5CqgHc24uCoxdBYOarLsHmSukX44/DuNtLz1qnOQ3eCCK6UTC9lEyd0kiMxJWlq+W+WxYF+I
kVeT5Cwl5mUIfIfdHSt00QURMHguj+s4E+jak22pBCFF2IAoLXh3CwXYsJtCr0zxMcQpF4v8dwFX
AgiliFpEWKPI4wJsgv/rmg/sYP62Fzh5ppaRrv0YLOWUDUfDdrgqGG89rrcN/QX5qXgHmvCPQH3s
Nk4Bz1fINPtH3YHj5VHGUTF65xaGjDkP9tqRgkSUZMsO3k92DC8s6y0U5HTovTH6lkCMPBz4D1ma
c8jgWf/eTLQUW6YpIoWUhFt6iY8TDkp2f+dhdnL7W2myBcfpAzrPrDa7kQsI1O1V8K2APm/LcsnM
MWnQnP/k3rSfnm7ffBmtowbAvpKSnAQ8fT90x/J0VFt1bAr6Rvn8iWrWlzB2FmlB22ucYtok8fZB
MyQixjbauFufOdgWBEeaST27ZzvYjQNMPM8iLxl8+Hvhowf94jb4k4nDEEQvBsi9/k86LgMN0e3c
mV8zQhSIdpaJdjGgYD2e0zYusP/X9GrTph7XN71cHC9LgOMjCcQw3pjweXm4ari2S3hwaHhCqcDt
ujmLU7wHpnZZ0FkgUI69psRZtHQY9lLR1htHQsVU54hXfDMvU2t0UQ5Kqg84TJuQhyNgbMLIS9sa
ze+seNm3Lr3Wli4xvwU3HBVuKWzOsLyX3ImZNov5M5fIe9/09NOOqVlbW7CyFrAXlrpWXAp+oFJk
3ZlThi0t4oMSHzjzhRcP8kXdh9FE74PmAAflOE7eYnSKDFuL6R+/YFZNeu+6uUNsFgrc299jkW/o
5r9dTRaialPLSE95UE4WN4QYXbXdGxnjVLSGfqc+w98++PaZLROBWPXcqjC6ir6OIHH20DS9vqLc
WLttwfb/MkA1lqOfIubauHxmO83PL567Teeo2h4JwyZe8qXj0Ulkz2HOQ62HdcLRPdnYD/7kXbAg
cK2GHRsjQhtm6jabQIMN4suidzhs0K/68QOOydF9ilbkF8BeekX84AV3OtQ5JSYvRppbgvdL+lLC
zXZwXLOxRz9R8dpK6SOmr1KDtCd9rn4TKeQmXzw+ncLjTFz6nc14sYUcMgJE0d6zjPWC3bF6fEnG
/MLhFDQES3OXinVsLbz9IYllgYq3eFFhzXCQ0B9XA+B2ByqWLdXy+rgSraXAU86dTZSZdcoYOAkp
XuyQ6C3IAwID4jw/jiPgdhWvIYFie7+jBTDfGOnuS4TAmSr9fIRDxXMu2kbAbyVg52r++/5+5LR9
dX2WlajplSidAzx9iozyK8XIfrjv1gSmpUDF2XfYy0h30/IHuGz95ZfeQgB1W3UBvUa/nTcQ9K+9
uKVc0PNJu2q6yg9hJB/gNOPNqENma3NF6SiAmky+Ttu6iKS9ELOwIo0QmuEpytAo+TycpQh2l/bU
9k6Bw9hMrN3bwOccVqzx7d9woWLZlSY9ZySE8tJJZNixXr0buLIA+3X6Olokur3QNxeM2lnOlLt2
e2xCCJsz+/C+vNOqaRUbVs1tDqzKILUhRCCXaEEAzSwbVcO+P3v+em2Q/dmUKMum9H1JJT+ktXr7
Df106WdXdCI5pDkE5HxrAodMTAsHl05xMXX1DW6onqsg3DHSM2ywWMdcjwiQ05LXJ8A+eW6/SbMG
lnm7L6cmfZJdu1LLCvGp/eAD25BsFjJw2ZLT3UbMarJ7I/Y6yr9zqZPScDIukbJEPz4RN6D95yqX
vmQesFfwQUoe8GwWIvVSiv72F8xs0U+4s4z8lVOb8AQiRp8A1zAhaP2+NItdSrJjC6/fwF8klr1w
AIgM4HlJkDaa2FTQRDCWMUsiDBLoEFcuFSUfz0dzr8Jg+XnbSGjeOSD+hCddslD28WZmlsFkqxZq
tVvHPhp5pYXFvbXIfDdVeJ6GSv+fLX/uilYetDCMlc4LUL8NMfLOuujbg26xLsEtLCJdv8zJI+uK
9wXlq/Dim4vbEYTHUf7pHl3pPPOiBMpz5pdmVnxXmVoOMjzhHC9TYFUa7bkbGLv1365dOBNRMP9P
adhiUw9+xvWGvVF0xof2SYhhRDUBjVCenzGI36Q+vpw6/SfJpz144gTcugF3QQ4KO6oghUl5Pria
4xMDxWe1xO5T2jIu0AKrA3U8WvZq6Fsuvaqrf5/94rSdCfHVZmvvFYemPs7uGDNE8pMAQDrAbTwR
u74yrDHqLevLlUk9r5QFy4//Y2ws6xtm8yREf4Gbp1ACLq1JVcwSPmQBwXGRfHA2vg2ElM9sJqbj
EiGe7rZIlRXCgA+oFZjHOVOW7fbKMP/fo8FZV8OzKqsGJTLusgOctH/Vl7gUtC3xMgX3yDtmVc5l
IX0KtOhmyMvaQhbtC7Sv4ZqC91F1WREz8FG+Wc+8BM84OWglquvXMEZc7FEWAq9dmPQoHuVXKWn3
LBcNRvgQDIAOX59rotGIp9ucCIhyaKTDMNwUI+/src3v3xVYuz2c0HMx8NxW3mNuclV5KLi/VA4d
xFnoon+fLG7Td8sSBMl9e80O5KpHz1akjnYqJmndyG9MIRgHC3NfCt5lfOOd/mCTBfotL540lqM0
m1WQuypaxHiCDz/yksDguARJHZs5lCUlYzvWE3Wo5cxtYLp9C5HiUFwPuFpQkyNADPkJQVgsOOyg
LwNhI97Xo3zdvkxXFFvL+371mgDv37ylxXdXI7gaFfZbQxPGn8zGTB53QzXEHFyooLzWARCslCvI
BRPX5XmlR0vueK9erRJcWFWGuPuu+Un7yVUOrUt9Nj07PFJTdvuBu1gVz/AM3JDBu9NJyocLlOzO
/0+UmfhD4FQCxRgzjcFdp+0u+gCAu7Z919r0eH34g3DseAtn439EaWn3cwinp42xH8rTIdMNhw7M
838t9Iq7HQPvDVpMn+dD7W8blhbsFnDSuUMIXJcOPOiIiDT5rRwFAIFMhIb8NfM0ttDofnddJ83f
jVxgtWlHw2ijZYP0t47psxJCO0dE0iebYoPw8YFdIsaJKTmMD9bcvqBAzqYe2lYK+vf6CWfkCwB7
Im1XUiKHddsxwhI4AXMfWlmV6ZIw3fga/XmsJAO7Hk4mH8xdTi2yrteseOT6VOuHARwJXu7oXhm4
Hrup+4tawoT6nLyMAeVemmiMXG3Krs/fdECRJ0YrzfHpDyXdRtNv0V6fSxehBZYju1wHSCXddolZ
b8gOjj/oKj0bUc67gyYGpQD9toFI+x5sNgt5GflOfy4jct2V64x0YJZTSpgWHpnbMQGx2sAc3x/W
FcArH9BGWh7SJDRXgFQ2DnnVhkcvN3DKCQJoinS/Ud/VYlV2Z5EXCMb2xjeCdWb8lpaR0alYmFgM
nnCyuyBvvXsKdr4QykeJ+6nzB909yaeHUAULm2cuBQX2Ee5/2HWKwbhQSvJugRDrvhGA1Cg0pJk1
Ap9ZISGMcey+LfIhS0s56IwQ6INkKAXICDJe0M6DCrMcISpCI/+q/f53RtjHNvcdxYfWV0uQvTje
9pBkU/h6ar666MkZJckM1m4jYWB/ROfYN1aMmfx2SDo0CRUIb33Aqx42/yy7k6TCyRIjM1up6RTX
fxXw+zhpyzdXeO3KuC43FL5d79jDUAz7Y5ijaUYdHWdkf3M6tK3wOVH4DlMLEQYaSNmK6K/nBrH4
8vW4I3Lrp0KXVTkqb/EPsUpPG5y243P23ZAepxhvOpXDDT6FmPeDRAN2R0ROHRQRX9RrTJlCRwe7
KJZW5bpVFtiYkOkUmhchD2QCBzu8sW5veeWnvevwoTmS3SgfuBqniGl4fGy6gjjXi8McgLe2H0CD
n6TEQqvVQwNFynj9TF9uo9OBp+bLYfGxrcb47a4ShxqV2ja6vKsg+XwKrG0lwOdjNvjVzJ5UXO62
I0eBOk8C51reIWqBdNsi/I9y9Y37gKtulKYeGgEKn+n+yfrQ3hkmE/Fxc0PyWQFUV1OVAwSmip3t
lRrwM4MLExTtYYSHhWQRlBK7XhJ3NgNgnQa5vdWiXq/VO6MbJK4nBVuoi5jWJlwSSSk0hvinK/X2
KseakAwCXbdAXXYL1Ij31O4GhwfoXA9ndiQdB7XH5NZDx49t5vBLkuAtkfTWmaYlUA4LCmlaWBDH
8BtCCfjGp3mIG+Tn/NE715Au/jjfokHFSbf5VQ5jXmEbKgjCzoyXT56QRDpApifZklhBDLSk7uG8
zvlo7jG8kuHYjTEyYMqprGTFjg68wl3lSAZx+Bw73dWIs8qOQp30KrZTypkN+7a4iaEWj4j9TPR2
NThS4n3cr2F5RXXJOMu7uER2qKt720JkUd6qtM7BGuyiLw4av8QEZjvjdcIcsvAGkwgGJWlFuFnz
MNGCbznqqFFmFxLYlkWn1BphQooiL4RutoUuteWKPnnxYzzEkRpdkYRJCsS/55EZSmoMrbMyMGBa
vKM1CCHOeKVaMY0krTamEzrPK81hZvF7I+KROT57viDT9qqO5iU/bxKwnhLGT/sILGq/ZI0GwgY9
K9G7kKTfSj/WUyx2ZcorLKjeTNXPyEFRolequ/Z/rLX1spaHRsfuABdVuQV0ksrZwH/qxxn62X2c
LA52TKeNULqZRLSZ6FU6j8Rh7XifimTZgAc6D7BAUssfjpg9+ktxx03xexULC08DxrB7z1jWeOjS
K+hzJsmg7+2baKDYtvxtW+4impfBUSDVAB4xuBi1WGSQ9tuW0uwtLzrgMIsfpfyzE+ZPuPRFgbSr
yCxVIO9qFMm8K4FPe/rQWSfY44QN0CHCRGH2AIvwLFJmGZZdsoHSMgmTvBMWVgVvha6anJERlgRs
FPh3c8lfNwTb1sCuwd7YLMbHTCrAxzpRgj1Lk/LSFSRBJtRvUjAyZqRYOlC/Xwz2CYHfepa+moRY
rn2u2bgpmYYduWSi3YIafmBuwvOp9yCv7X0DnTIBm045NQwIarm9MpUElawkRa2dsaFdM0rM5uV+
pB2FzXxH6m2T7lyUFQG0BRBY1nFx2a4vRxg2sz/JYoSIJfD+VNGyCEH8Y3FipURvYDvKPUDUQa7Q
jD+SflEXSc7P5q+j0DtY0mMYnamqZmaOwcMHdtX5vjAECxj81TWgMANwYX5K6a5izxgEFPw4eQaU
Z0rTIYEPoTk+9So4JGq4i60z442v4phLoo5sMv1M7XfeM4m4S6bJZY44X/TxvhvrKzCZtty0aGvP
RrixezCgeoAUxmJA9YKI+WkjzQwxaZyYFI4OPByS0uN401FanR3eBKWTELCsXZxUB9MJ0cVHiQib
CoEy3pV0/FCLhxfr4dLN0k1DC8ET5q7S1GtR7AVyn2+Mezi+iS8DH0Dn+Yp7tfq2EjMIddjmsfh3
I4bz0db7g5KfAK6CAMRooLAvpnVDu8/E7QJ5I9VWzsiEr6PC8LW67CaMlXGtnN9azz+tKbZS0U+O
zvl0+LD+tzmk3f79JOZ8W6RfF1V9FASiannXVn3GzrW9MN5eT1BipjfSgZhMuVOKVQOlAMck/kZT
xaNiqeq57bzHu3YUcV7Evz8+LppcZY3ZLRKPwoY52UwqBuumDQC61Zj85jnVj1rtr8mmRm3WRmeY
dwwZXnBUvvzgZ5z/qMAEPdhhuzpwxZvk9O/peq7fju6PAOv83vek90jUvJychQj0rE3InCw0uiTY
pgDq6//JRxRwTVczljevoWYY1qJhDhUzR1osJY23cHm8gAe2RcIoAGyvQ0bAGntaLXENiWWkcwDT
TnddvqkRN+wKaaOk9ZxC5Di/5UKmXCanaKmuc+GldUMi5nl8Z+eprO7yBfU7vXOmNmq5TbRgVFvr
vToYzrAVObTUxgGuECMSCtkHHAYHZdWg1jsef11B+jk6bka5+EJ3N6slBXSVcH9NyZ1pjGOEImfd
mqgHJ2oJJjLVV5ARFJI2f+gbihNJgceR0ad/TipL/YO7867Az+nDWTm2elM+mhE2XSNLdvgFAmOh
bu78NHfY8tTBeM2hCW0AEkpSMZMyZHeNeM9n09vNwvzwneh1V/EJFtj8PalbVhduI24p5NyLOZKt
+Oj22cuqm69Y7FpjJWAupkAbhXH3hKdRQx7v7zn1ZkWu7GqdOOfGYUgmMCOXOtGu7c+VDoMdKYYG
4XAB4gEjDXb7daNmoSZNecOTLqoOY4ZWZWIMDOLjpwSvvYNDizKQxPfgmCKVIABvHlbS+2ELxHwW
MXruqDjPDyAFYB83Q+4ek73GACW/5UawbIERZpqI4HbiXrybt0W3FMgxKpkrnJHwQju8NsFqgJtB
SeJODB47N9FV0TfD7VpJJSRHvWoyH0Fn9DDNFk4K3KXjb5XQ5sgDgjBsp29pdP6qcAX4Oa2Il1zd
3RJl2shdjZ+Ynn4wGOxFxbC0uzVMADyLNHh7i3ErZWDpcycu8wgUwOypCxAUEzClmNl6h7liT7SJ
oK+Y7kIuUnJybj6uW7z5OQObML85UxclkYR28qghgECS7DoSYGAL1NAvf63a3Qt3txWK61h5z98Y
IJUsfW0wVn28LgiqUM8G/BA44SWAz6DvfKWeDcjRygmD2W3n8TZEeexV1Sr/tGSnBvwzQBMnL9BC
EaT+Qs3TKGvyw6mnS08FVa9Aaj1OXcMruccdEY+EpAUS8YIBZlIYK+egx9a7XugRiQVZngvSrzYf
VGmAqrljQEw94a+KXE6XCqVQ2mZxU5jAYmb+nV/y3nCyupvotEFRikmNm68vKpjh5f1sWX3/xBf1
SPUHcqrg8hqfiWH4w62Eumw0oFjHYqN5ZbDy+LFTyxCLRLu3wHFlhgOQfZ9cxIbWT97lfRbCHDoq
EJmj5r/5B5PjeWjHi9G8VdnhiAMIvBw7wD0zVhXlPmGTLI1jnSQ+LZ9qAyZiWLes4W7S/WkVdDA1
KYGfD0jSyvQpawNFi3TkL1cL3gzHU1/5NsZkFbGbr9AXPKX+dUS5597O+CuKeQQc6EzZh6nqffwu
JSzNUND6A2RmgNeyQnnjGiRgpk0Jh+Hcc3QTuselo4TvC/SSt9NfoSWO9/qpHktuPmubmMrQGyGv
tAQWgnuOiEBov/YysThyts37lA4trgeY1s8Q107Dtt1n6vXxVfHfvxTQ5Kh9zqighg5BdA8lAaEi
q35lhMukvvz0JKwgx58HiHg2gzoMz/bSp023TyLpStntEerLFxmH2CD5lpGfXgZia0+neJi3t91B
5PqteUQ//QHcccXG2n2pYip7g5d5SV29MjZ5CH3/2zfqTajKp2JKmqpOjCg6/oihQdaEUJdnr/j+
M3h08SKS+qgeF9ce1ySYDyOrvpD0ISVFFIzOHpqh790igY3uxTqaB3i+DFEHcLnCMwzcCmEjS5/a
0zPVzWn43UObzzIv1hOqje0dCebVpZL3Y2KeYR7Ki/ZGn8poe+//0HdTbUK8Wb2BBYsNnKTPyQEp
POCCFuv3J2FyS5Yumd2Yr+FUtCqLBHY80XXu4fCtOaE2u0afOD3rKQZoe1vG0eFRYG1CodC1lhDH
ikQR13f0wqXoSkkm0aRo6ld3WOUdD4KR0eTfBWkKdsdaGoCktTYoihOQUSDogHr85P3mWyHcg2ls
OMSoRsLhVV6Txf6nuSU1/vlXvjlTDkQCu04+M6AGCqjqU8oPyL0/y8urUkfq3nygfCYgqWtFZfv9
zoR+BNGCFznZPGO4dzjIUluqsSNMxeJtuBe/rTwsCp0mUJFkKx/Y3Sf5P7j/2vvBKuBQKubrLzNO
Nom4g6yO1vErWXtrSeJvEJAqJKz0+sozHRqSubK2FJQxHY349PARN/vw3Fhn/GtqOnSW93CUTeU8
9oE87JxUioaQ9e1b9iyO8VnLBu7GTfkFbfQOxMm4cTH6R5RY6oxbdhAkh8ifjsoQT1X+zXKzOu/j
2xFwBlA53wFPX0lYkG6+NbC71sBTd8mWOErpWtrb+AnellaxnsCWgM/bjl0RMdRVdVHxYCed2qx4
cNHTqtrk4sIJV6X4UblfLzrkgDnF6MMGXh8txxKywZI5pluH+K9hQMlXZrsfi3LjNCXdkrV0E1xj
zyXrY6f/Yemzf+r1nxd/IGAbf8dL9Q3OQ7e+lAFvOl5NKYzpdQBQoii6wAcHmPv3LRSZ0PunjsC4
gFhUPwJwCc9DCunIbk8ELAK9SkpCjf7WaQRo+Wt3nDphXNhnZdTBApfQF/0yiuxFaOGL+nHd0vAH
1DjQTA0+4VlC5K4Mb5caG3rTftEZSAjDdCv9OJkgAU9dAGjESTmJjAAA3wh0cltKf8w8VoNHdmto
+0XVrph5o6JVtKdBXzV0KJk2b04bIBCWnY1DwHR5PSROKBsvlTcgaGhhpjkO2tLyOjTA2bL/uY21
Gy2ygL8piF7dDOYTh9eOn9X73Oh6+06f7zBa6VJ9F6VNHDoZjuIsc2B0FZJwWW4b5Mt+BUIAOQls
Qffgvx9CQ17Hf73kueyAmgtauA2Sc33ekTEM5zEyVxGSrFNjyBPssAp/07QHonBiSWAiIiwgpsk+
HG/dK4ewAwjDlzEdz7iLCZW+Gc8zQRpe/Fdx+oA2rpCWpZkpio7mT8zJm4AmxzYKzeTrxOl5C18K
XleyCX6ipTlfu3Wzfa0dsP34I3nMaw0pDH63KXxrLzaJ8bUX3VeY3e6PcVCZ/cJa7W/4fj175Fr9
I2ZYXywWd789UCygoYArymKFNuaQ6M7zZHeqiS2ckneGhp/zbZggOkOnDsmTmRnwvx5TrmK+rqP7
Btv57jawxAlA1b9J1Lc1mtqHUB2jnWkLH6xAnJ1JXlO0jOLxptKcnXJYL/0Bynd4NVNosO5fxB7i
4YcpVHFTMrtZMKj4Ugjy01Qn1ebneer3n9mTpipt8pyC/ZlTR6iA9i5dKFuAgqtP6zWwBhAeONw5
zAjlF7EBdCbvJZvRuJlmGqUdUU/6yIMjRG2C3VZ6vq2DRbkycEPrI6PlWIPgo34hOfgm/pnIlWu8
MsA4b/m1DCA/BHlN5B81PYZ/uta8OzAVRsUEA/0cVyiI7OAH7CkWkpfpXP5WdkZD+DPIhvDOhJtG
7teA4i3/3Q/VBjlr5y1HAtSxix0OBQPFH769lG8ABkjlIBc7IKv+/XFmzEn+LAdXBdp9kOPkamWE
rqr98krjZIxLrxgrN00aROXXUUbhqxpRlnDm+M5BECWdDjaf8qF6QVWc9NgcQh4XZHcSaA0MC093
AbDyut0GqVcADECKIgHiIIGlfNKbFfxZHwzm0doTJ7/7y7+J5TABcn2l1lyewLWPFQzr9ZfshauN
pWtJ1JBQtKfnbGx+MwQehFOALAWeiY6FmR83Sy4WMQfqIGoqP/Nc8ALQJ0vhu2YBfUVdxEXlLwJd
rLNkhni8uLs/DGzW3KttmSww8NcbYd4BCMAEWoA8J0utZNSEeJg23Va0gWpLOEJdjsKC9B9UMBb4
ztgk2DCtJZLiDqTc2f/3+nXW/SASAPiIWcBk7hTYK5/slwfzVWszrV4oCZYHIV0acmF6mYq3HxMv
/4DyJwQOk00DJ+rrDONxlfG8p0YOh18+FvVxvNhCeYHkinm/VNuTz0/q2jZzZh26HDVkVqggKa+w
JvOscJifJQpU+nmiBpm9N2DWdkhi5/TrwgyFS4T8RrA0IoUYXdJSifjVyd6fIjyKcFZYPmms/yML
VnK7Om6evzq12vBMrhvOqnlVy863iWafW2As1hmpKaHAr0Vs+zBswA/KR/k3XFmDl6fEV0/mx83+
zFx7SSCwPYHE0OHYZu/J8wUklBL07erBeFneC60ll3VCznnZ1qdf5hvtq1xAO68JE+7U0p/pzX+T
shQov04m6chO0omZYrADjCmLE3Jc4IMDPFMYdSnW/bWyQrEUwb+8W6VBy731xthBvUbFfbqOv6j7
4MBTAfaqdd03zW73YtexFRQL0MViEUDlMOaAXFBMSqGMQtdhqPsL8L5Zr9Cl9Smw8k3bE3bwDbcD
yf8JET2k7qFdOCKmbJmSothXwSIZZg/40w6IBP7WZ8fb468D6NCCvOOjocNEIfOqU52l2+hsb6fz
Pv76e4G/qkuktBA4sDckKOErHdMhU62mtjNEn79G6Rg9e5tGi4NRE0ihCr4k6r7A++OxTyyQNL0O
J3s8i90M5RM/8HYBbmGtj6m7Pt8zUjTSw+mZ5vN6ToDRwBBdVoi1wObZZPSJz7NpvwJDo2tZhsgt
gruQRHfTVGMPqABWfhvMmXs4YDPKTXmvMqgh78dffGDWm3J/aiBicdbYicw7omaljDBpAdOlCwR/
nvu8AnjVKkUJ0S66lSOaUto4q85YWWnb6wgGGRSzdXdJuW2abbgZ+cvCI9U3NVI2gx4gzDg/QVlt
lisMEtJR7OZVAc5n/u39+6oFlhr+rTwJYv5b7ITwm1I00vVislCVNyKpPZWJ2INZLqgXGzbPK7QV
ChLpRMTgkWjxOwzdfR5Bq65MUUmdt5yhQ+aAFLrxvbx2BE6Guq671NdlcOl7Hpg9Fvlq+QsOrc0f
din6+1KqVNG1tA3kiNuJVIDFdWUvsSxAwp2k+VmSkvLimrcDJthReS02M8vwfTzx9hAoof3Gtqqq
WxgrrDDcjQwkUUxNHxa8AaTG//LTxE6weW2WveOvQS3ylY4GHd9Y3KCFVm1cRa1Z5t/FcYWldqub
zMj1dGvxRURI/0W/42oWbxlfLIv4JW4yqwmRzTnfJuHdF28R2fINBVBi5I/6R0HOe16a6L1AIvHH
FSDUaNGeKVNQedN1xukn5J/tjgrLnnjHsvuKBp/YxtNXANOs89yi1Efh0tD9Vh2N48d18SFKVfsD
H1k7IdxRhDP31f/r6zUdltPmXO7TUH5xw22b9qMwJ7ysBPgH3R9GKLZ2lY3xNb9ai0RNp2Nr5Pp3
rnDo6GTiFzeolHFERaN6MbxGDCl5/fxdgXNn2ouGiYbq4dinXmqCToCeEWD9wl5jhOsP7zBe3OI5
eSf+prquSIc9MvgG+9UaWOrGAHCJsU+Mm/LIBO4IlJSTkJ8XOe2E8tTnlFgN4bozOiSDUSgm2Kov
is9neesmY66RiplD124vTY+Saa6DT4U8jmP/UWc7R5gRRvrc1IvUNJLPHExbizAfceOHDghan5OM
PqpGTItfQeNwpxEmmh+ZAvmmeGfkhRF2da0cHPfzBuz+s72t1w40xk/26sAknJ2t6ZdxoFUlBhS4
SQ5AQYtneU93bGK/EVUQEebLD9q2ADDoo5M+jJJxgNub+YNf5KL+H3SGBvroxTPfcGUefFtN4lZG
kW6UZobbk0VzEShDGYbw+/zov876H25bTtZB3haZ1xchiMvljN1cXTzpmN1kZErGu5lxzsBYknv5
4S5aJ2qURNPEQARzF940LZnS5G4hM/XMhQjzf8Js5ap5sv4amalYg4aoT0vbqxKR9Mnle4LXaD7y
7JknO6dHRf/O3gRXJJaUmHANIhlaFJze/i6iinv1hyPQ7neC6l3+Sboc8pWMheB1G43d7bJ8mZfW
OGxSoy2AIHGRZEH7D91AsU8RrFc81/eXX2AqYhYubNVP0fm8Ge8ovuM6jyBKnVI/V2HW1e29uoRA
NvIz9QeaC1KXH446WEH9VDbypPpU7rgqFrj5VwjOHoRjlk5gqfu11KDDb4uKM+sdV1yC7nv6A2jp
2bY7keFpTIENXxa730r1pJ9mb35T6Nq3SVWYRAUls3+nAcdh3yCHOdiDGtApKZjbOfAWCwb3gHfZ
85qDBDHpcYDZImEl9asj2aho3tXatvnjoIjrINpLY3/1L7YNn8CQukL5EsNyHWL0G1iniPE5dG8z
Gy4vGLup7OOnlE4CwFLDL+MSmFx0xXqu3Uqa3WDPlsKr+MFEOwDWZitsq+Hd2QDnOJBmIjUy+ter
A/M6ugaSiCDTpip7+7fwCaqcvotTNeKQj0Fp5dqn7IEdcLkpGavGELb2P7Wk6o9kMCRFlK47kvWD
jrwbAkM8GvSoD11SWf6pIKeY3umyeBqH/Zqfb7lo1gUIKeFx83Ph1y23DdmEQmYyd824unVPmVTi
/TwEp3ChX7M84G+MFD5UsXN8e7pwNwNxoRw/N+KfQigIUkfiDarPUCmaLuT/U9z3QkfnEzQYI8P3
YJdjMaMeo8qbEjS+2EDDsX5UupL8Py4LO3oBriw90ih3FjjMDOcc+3aglZOziHYSkD2V6ff3RKZM
FDvzCuOAEAXoqps5VpFxGQp0ofG+muNbhEKz+kdb9xwqHD6spz4gKlk5LD/FU5iC9RMP91H6RjSM
nm6GZQh5vzJw9ZIf2EOrmPRxKBxkT8QBkClr7wgqKJMCtFYrNX1S290sVVNUl/lobVUAblDBIT1a
yHi4xkZOa+fqpTPMNTO5S4YNAOleSFYvCFCIrOlU1hTY47KmQ1eEfK0s9f+bmW8hbmNxJBTAAgOX
3+bnG0cm/CFgzwbsA3AcQykH5WID5D3TkS/OLlFLyY8l57wL5tWy+qlx+59iEtmqqjoebqdbS1qw
6DlYVZM1S9k5MKTjrHtluAYgUMoPcna7gkkYqYFg/E6K5OeZ2rbRniPJQ344mBgejdONxn0oTK4j
aZkxVNueF/lM/7l7Ypv9QN4x1Wuns7ZJzQ9ko6HiDo183ALPz2lN5CVEFDkOzFvyladEMHcSdZjh
/DArPkDe7g2ibznASjEjmloLFmbv4ZhvbLt9x7eiD84D4Dw32Fm5V4jVXjOp7MEDHka7w3Hy484V
3CAQA0hOA/gab4IwKMi9m4RPiITHQVmDgPFeoi/HdXzS02uHcSDUmjewGSGbWuHMsoWJ9hUeZ9TM
/8qOBCESL6AE9kR90rTjI1JD6iyVWkfMo4YzXy4MEa6f8fNMbUJCM+p3jZZ4aRlNPmnTtH+kkrHJ
WA74Qjwd0LgGCScPqM67C6cUijddOhaKv33qEn28wBspRY1njrj6Vy9Em5bHtl9MjMQeQWTeBCvT
HNrlY98/yA1EPrZ4No2CeU9trqxCeGim4XeaoERcsVsAeQLwRFrVn65S1O3a0/8eM/ilZosxY8CG
IuKPn9AUAMsrmUvaopzZ/OVZBEY9LcbY6bCXntXT0pwRBDGR1H3lF19elq7jYfVyNEBhAT0+bXs2
2XYOqnQJaDUYGO/uCrGwjf3vTFbMr58Pams86GP1//+Y1DUBAKAXyjB9cW9zWs8WbLmGRTJAUB77
rUr3ive2GSTShXJ307OEk86lYnb63LrgZdRFObP8U1l7TbXaYoluB3r/druxylHY+02tNLnMX2WR
hMMYFB5pxcbG5aLWFkJCXiCP4KsSjiEgW7Uz6IaJKMq9aTbPKLk6z8KowRI6a7IYObCXdvj8yOja
DKMTL/A3BEiOX8OvDZlnziwLSSAGVVUJnfLgkr6XI3lhSlthbRNj4+UgzL03rgo8hEBxpvdqf29M
dM6zYOhoniK1TcZbdSpN8/QFEL5P+ZBi42Ryt1BQS8FMRW3/wj+lN1/9qsT/JmNHRT5Ds1yr7L8c
QeMa5uazshUP76ytJu7oMtExIT11fVM6f+34xCEy0U1wouHlD1P05YeSN9KDJnVR24As1Gaqn8GA
EAjkTarlns4c9unxn/Un6+A9TVfHfCrNlTFhlO4yFtbFPSNNDStQ30i8JEjHCUI1hZQJh0Zx0clW
XQa6fdaLKjD7sJg9X6/eTkimoxwDK/0ae9oqVPmzpnY7Tp7G00yEZ0wpfHJbCoRPD55Pr0VT8Gj+
p9FKqpOKsB8Z1uS/6/Cee3JjETQWszgKSS60QCN/Yrjs8RAi8l9x5arh3N6Ml32E356DHYwWv2B4
Y67DgGRNLFqkVJtViVU+U5j9OzKGsk9+PTGsd3qSc6SSdBT0OUyc9j+q/OZnApMuJ9Xt2TI8XTes
jxULrtIqr+UMDPE0H05Dz5dz40wGKQy9CYemNz5e00seix97d6l4unJ+ig7qg8y9ILbNFEhzV73l
Cy0zs8nrGZDpSZOMSPI7eWz8D3UQeeGeP+AGrRSaGGgeVlkuTsZJDnBJbm7IElXfIVeOvf9IjHcW
QBxGIt6QuUuPkfROjMihSz/pxSqOmnCtj4cNb6DIv0so8oLQTU6FZzekF8pSA9vuV0uZClClanzZ
Fj9fErBTIisDJ7tpFDrhyqA+B+wzlruyVCPKVKQPX8cXVmwn9A2Yvws4gILwqPJsugKaN2nwOVlR
hRtIA5osh9TN7YGbjGPVhV89DE6Jaf6QCD9wePIeDAWpyD4jFq9GuXHMU9rupW1rjryWHmHCdeiG
gcO8itJo/RmDers6tagWDs++TQIFc8iVNRJYlTp5UxbM+qkFjv7/7+b/SX5L/mb7D8bU4dlnJswq
yWNwUPFTOjSg5dbqIkM+g5aPvhWEXn64MzF+CY+wcDtnzdPCtGh1atFyiGtMfStFDZBuaDDQmuRT
fnEhG/1LeQJhThSUvkXh1/7Gb1gzxGEUgfp9+zddByhYUQX0iZO94kJ91sdSgCTyOxYL6Tg9j3n2
o0JGkU1cxS3yBI/W9v9kNXRmVoy49I2OsrUcrLjBQAXedQ2yOhwGlSyzL+eHMrgUl118reRH4W2y
LBtdXBFAw8ufVM8Yn0fFr0xj5T01d2c6nT9ucbcWNUAIYV2QdqL7kBxugLfx+PWeQuKcZg9UJwNW
JMh2yYHyUnnqdoITtYvyyeWQ/qJINt+sKeJAVVPJyEQmK8vm2EAENZXZzU5nkBNmmfWRD5uXSAwb
ANvC5f4Dn6VX3spYBS6tLILw4NbFZIWB9WyPQ+oUs89WankBYCsxJaTJbWTMBguzA4dJo6oMoGfG
rQ4fjJk9hk9Aj59ksq71iYNHt1HmlzNKLtwa7TFiKPaKIYj728pFiaycTOCex7gcLHOIqxy6DKUx
bZ6qY08y4Fp+LmzYv41o723wvm/GJRkpz2fT5MRomCmXroVTZ3Mc35fGPHLdajVr0cjLGOqov700
ZPHE6qqm+XJ82rQnMRfhFcpf0VamA0IKy3Wc9F+lna5eFHBO4axIQuT5SOX2BTL/fpCWapsQpvKS
99EFYIMYQBrHVVHcWA9kBak59UYEqkQERPw/fspQu6CB7e8+HakLCMoCPq1bWGGP7TrEsv7sJFDP
zNNHcZJfJb7Yq3OM482OJo0+JA4FpjTCMPHtcKzHfrs61D1KvuzvjUhwu6Tppj1umjjUSh6da5ey
/Am6H5Gzq2jse+Ypwdl5+be0T6+yuupb6Nkifg96O6VXiea6yED2lhYgdscEk8yyfb3Gvo1yxWR7
S5bUoYQh1qvZ9dop3PvYCfVntQyJ+vjLzeL2pl4xWtA9Yktnsc5TGZ9zHWnf6tmrTEM81A42IWFV
Xt8ttqsOwug1erLJH34zeVJZNTIQ7xk1bZOl0lVRqnFHzbbmGu3p42k4Ejc7QBxZE1yH2+wjmvPQ
w/DFkW3D2/eQUDg3vKtvUgCCTO861RocwTg0RUy9DDOZtn7cp6nPsEF5G3C0ZeiVVBEuAvDzFiRK
SPv3/vJ7XiTw0jJNuT9XcH8KzeqZi35gBk7act3oA7VCQCzlv9HlaqBXW0WYxV5Tf6Bx0n8n+PKC
Papj8Ery+5iSKoC3fhDabk7gFGKtUdp/BQL3q6JdRmFJJaUNOOX2onM7rlc9LG17c6oIFV2qNYRb
q86u+Xxm/e7tntQNiJD5kBT8QRwG52jHSmkPS5Dql5IiN4Xmj8Wpbh1fumb4GzOn2PI41TTqbNFk
UGdkIAaEcyNND2KICotbtLbioZENyduUqkVemmhDw+sI+KbOQOpwQ1+Eph1xIlMFkeJGNEER7w/R
eVl4PLkfldMUvw5mAp/GEVoIDynK3BPzzG71Ro8zWT/wC1NjG0R51i0qOzOTsbQxGvYq5k49IVua
87WN7o16qyvPjbNONsZXFm8kXNT0Jgq555LzRxL8Lm261icpVTIkRbIZaC9WeJ0nBp9d69fXgtmY
ntFw1E8fPuJkRwhyf/m57JBuP/37GDrXQLoE0G2qHFc7GTzbgb4ZsTgv5ishKBjSd64FsdlhmtDG
ESbgpv1phZvyEFwDykFXyEjxwLRuCgE3KotaKLwFwRXNG74L/CsYGC0SmIqQroPyVpR3nlT7ekCQ
0V+Y/QRdcNAt7bBayUc6oJFAngp0chAOfPUWHD1y958q+A6v4Kx9cILmFCi/1YPsVQXOMSzylH2K
RpVy3Xfjla1dqAIaSBAJfswv5taEjBurr7DXr2KOvbghwIj8tkgfGIXeugiPlxD6ZTAatBaIM1Di
XvJ0iu4CCMS0FIBWBQDcXy71l1dSL59Li8SjIy6Y6rmH8qAndGOcJ41yU0lLkSETIlRa6rErGme6
R6PEe9CR9oqynE2JvIPTMk6IEneRc0X2+2+0ZrU+ks8OoUH1tPgEF6mhyapkX86LYTnMztpe9ktJ
unr0ryG3FDRhvGy1eiuz6c4P2miINTIxWssAhAeIuPNAltGI6Srtm+1K1cBY0NQIqjplVyCiZFf6
03uhRivuj9HdtTeMdkubjM2DdKCAmcQyOdTi+YZ94oex+JHX+EmzbUwWSzzmiqEwwnmSRNIPu842
MaatatGoCkUK2Q1HIk1b5vSJZvw9lNrP20ndiqMSvJlTy8/davr7QbVSjsNiifLRxIPVoM1ZK9D0
f1B7AjPAfh47BICqqRpS0yTIWFndgl4oS/1sEVM2pb6dEu01dtLz/6bd9sNsiHVmCn/fy7HGPequ
CmQQcPz3KZ2zSsQSKkXh8Cs9ibx0oAyW7YwyK1XKo8xG9ITvEULJ0bjxeSM/8w/yYWdW6dKh8dn1
/qifygzf7oqI6vstDgKf7VSj3owLhaaSu/C8rTWwUQ5kX6kplLg7EBhI59AojYLzgdewcdOekuEE
UC5e7iJQUTPks5uhhYHoDqM0mI6yqVFeSLeBuHl0fOunxtFi28IWLb1KioCgtWw3/QID80qbL1SJ
CrTIOJrW0I0uCQoASKM7YHDyFtrOewBtkMWxkwSgovAXjVnZikYdwJsYeizsgBX5ToKxOHj4Xcne
V3aADapLsgobZTaUObLKDSVvZjqYkCbrsPkAQB+g0rYeTzuNk2/vxkO6hFPjci9J+H2dcCJ9MLXD
qg3TIC9fimnDkjBTC55c6IyblSiHzvtRHck6vfX18uYNs/WJdsKlhDZzDwInxRMaEJFjLnXtNzDp
v+X+0SBAz7VH0PDgCxSUKSg0t4jZ7a2tsddLvjymMQsiBYEckq+9dXC9j/fDfRH1OmJVSAxxn5fk
jL7Nyi6X4XgFIfXdMDwJReKjEceQBtTZPENhdjeLGZsb5YZh70/SRx66lifmBcqacewKhANL8bll
4yrUEMTc2tKqv0AIsBRvXmaNBX+yXFUDbxFMdJMHAqYHagQJDS62Y4K+LdSqjNlVZxgqT3SRjeFF
/O7MoEUMnLxVJmox7azY6lU+0LxkD5CLvRy8a0MKYH3Xz9bwWKRo9xjmVBMk8OVptLlwY4S3lb7+
NLe3EXXhO8Vfh1zwmyw314/i3wUOH0joP208b1Tw/Rsw2KzANuNYYzvByP67S3p2Ae6FN9AW218S
AONQzgaonvDB7N9dzN9Ea+TTUHiEPX5jyXAISHlQsdL7qi95Cgt4wkfRMlz+RjVtWBp9v2pBrcIx
utVnPtpWde+PhJNEK0IWcuByeRNUqby2hUIfGGLMZSLFSBEUtOG+WDKMd7kfo/ForlkufDtd5vZJ
vPO7j1jYwHiq96L3LZNOWE1M9AFEzv6XFLMmToDPtqDZVVZaUHrgaJdgZjv9jo8oiewSmFpZkeQi
j8O3JeIyknEUpom8TxuxcEx7Cf0mDia81OkGz9EtKxrPVkHUiVYrs9LEp+9RqEOjO3RSHqIvR8ND
GS/scID4HYqvrCM6d+CKIqKOeW6Mq7HlV7cdkFc/mK77JhMDoGzWNrPL3vUAKYFPLRnORzCLtERq
gTZAiIgek+445fIjW5gEmSmdL7iggYuctKaPUVl7y4bFuYXKY/Aj0hIatEKtywJyyAJUoTqobH6I
HJhZI43Mz7UlKtn39ExNdrASU6TJwUfghrQf1KS3u8N1aSTK/6cRVbI6zSoPxawqMtuF3tw0YR2r
/hPJly1PjW3g7IqEctIkE25hNllfnqZyeMEzrQdkaxZHchkQvyz8uFyFx98uQOgSiieFCH+23gCc
mDACbykFu6SWhivZCN3m4mK1PFtVOuxZJ8GuuipniKafLMupWHGsf/FtDQ9j0DW2BnfbX9G+jUyr
lqAn8GM80DQv7eylOuI+ut6lPNPemjZrIdQsWUUCY9HVZ1bxDKXjXuZVAdHBFglvaJ4k9ZwfCNow
aG4Wlnrbjm2SDebVmi5rCJE0ofVnfNG4ecVRYTQqXUT2qLb8aT7OTA9ajPJjXfqb1kkj5AhWqqDi
jq9V7/hdihFNVtJsRpwL3aAYCs8XNj26MNPzKqcPEokDRmDwJcRx30JleAGgXtjbMV3OBqpFad57
0dW3E/9FEgigI955LAJebsQ2+kRLqNojsqSCfJXagPboyYQ1VbYShoweo5OMKhSHP3Wgv+G09Kzx
qnK3j3V6vMtppM3nMidZxh42L3cuh7Mf4gYGhcqUr/f/4O8uHwdm/fNBtxJqWWcHeopjbRgIyutb
zGCtzkFf6iCKd1trbalExpGdetfkkTMJ5iv8fy6zIIWix2tUdiU0zs6n51RpKTWbc9/dC6PAh7GH
uc52dZry94inkCt6dsJO+69ZzkYlrf3CDH9sLFOH4KtDcXAKeGuAyuV/bt56S4V3XmWYcp1OV66y
vsq/1p3Q8Ik9RJiKyud8hL14BMPiY4y33oLQh+CUux9zZphYf1hS7ef42IXbp2nhy14HHyfjzPlS
QtRnOZjTJU8MywOF4JXb3FzMKe12EZpP9zFS6DynoHGZCyij1KElmHzv6U6xi6hfpz+KqZ+bdImF
XSEhUUDbPhF+KncUe+YF3UZTc6rUi0K1GvGwx44z+S+SoGyWSDvCydc+Po0CFbVxBE53Eeo25P80
DZ7/SqOAGkXHBtPUX22t3sg36WbZBexDCnc1/UHt8g3g07HHPZKVRk42j+uypKn29olAhUwR7dGG
/SPZ8n2vE8zIk0YL75wyZuy14dyB/vpp4+/0JFPsLCzQMDdO3dv6Q1+X0h+R/ghY20jxf8phZQtE
fEEZayLYdBeQ2pKTZNNl6upBvnmOThvwKvv0ZupJSlVQFteu/8tVt/3izsUbhiLItPFwQNqn1++6
FCRzlLpI4+BpqjPJH2zmqq3rJV58c7lyFjxm8cJ+Sjsw5GUc6ARj1FTLpR6Vc2u8iWtbWJutp9HJ
DFVVZavVJNCvzZblmy49DOq3iM34ziMji5iQLpDGbDAFrF5sv9sMf/kXZ6FFu8oFmRzHvO9FMMsy
SiwRIjML9StP9gtkgGTqb8LTqsDOQGv/XQwXvCWiVnYUcRyfYz2L90Af7n0lkQ6hyFJFvlRT8aGY
t5OHHlHE95YrVV4OIL5Mh9xP6/G+gt5CrDeVsZhFFk7NEeU+Fu0deNcMe3C05FmG/zzP0QcCgzKQ
X8qIBeYXy9/Nc7u70/VphqT+KvwHFqaxzV7tRg6dkNnHuaEpMiDCUQlMP5+uXhbONeu3lkbP4hnj
BUM92gresTeitJ3z3EvVlu456LpqHBiE6eOjSqoygq10ckbmHewXWtUF6wvS4kZeVm/cAWkwPUvA
s6lUDU/mJINZ6b/kR5a+9qP8rCHdrlH4iElCiuf1z1YtEQRvb2Jq7TUEthl1SN0ejpEe06jMQG1D
OYG/aSeRZQt3ExcZCf2QyNE46uEZzJsNu2ONoKxcWQc9QDwOkilal61pqQf4fPb/EWIMbdHNdIlh
K2rmPQWHy8WFlA/pJ1c1IjVTbBgfIp4IzkaQZK3zpgaIg44ig/N1tsu0YJOvbGP9/FKlBHsyGfpa
So/U70UmI5zy5Xql0WFv2QxRRG46CWSC+QhwpDSRzCSudRHBkYPDx2/WNXdWPacl9WNUVt3Qolux
zrw8bAm7vL+38yRvazn9hQW/2FQjcO660azU5EyAU1Cp03vdyp54Ln6DF2gMIU4g9Era4Hq3LGXN
HElnz72yKD2v/fdhjGt9y8oLikEzCQ+vEQhMTMrq2BSHDw+YhPrDlVnTG9FGG6dGdKIoasJsU4z9
RCnnPY8N1LEnJxXIUH1xR6+N19lWCRKp9eKT8i1oaP8OfCREKHXfTia0FYJVEcxV6ORAl8gymfhm
2nemNIh2djHzpENvD57uv0Pk0UuCLxHxWuHZ1V6ZD7QV1m6/t+4pMvc7CMAVq3OSFGbhZNjQZaLa
JKKjezSonMlds+G3s8ioBwVcAnWvZwKyIy6xhtPr+8sMdUmrSONyYUjxa8PHe06mJ7dx1eWP9K73
BIh+PbyS3zYIh2tnzBne87iix19WOz3MTpseYcaHWpWvAODfbd0GbdbViq/tVZ7yxJoKHeGZ5ys+
fyjIqAsTD7OHrnuzm+Y2uzvtCvywzO10rFHYMsmXjwXr4GtvxrNX/PGdPm2xbCaIQVRYhMHUNyTV
M2Wv4yt5+l+Cad0DgOzuiCmpS3ULe0xZ6AbIJiEMy+eWpVj84MX6ENp0aTe64PmyIvnQ7EI6X/c7
UfsGwwxf4fbkWlPj93buWcLFa02z48ZMXhV6w5RJAi2Tymn/GQZN+8EdqbZHJXvxkEjHbqWs+q6y
exzIQ+LK6w7jhy51HAdp2uxhDEsDrzNVnJb8UnTgHovRlf2fGCU1zKRqtM7gF/8JCaSeSPwSvzLp
1LTng9SZWZmmKYv4fZcfxefq//jh+kdq7p+Na+DTSa8abLctN+2L5JQdtATptpadw8DZfxxS99Y+
A6VcfrG2GVdP3L9eQLW5odJGqF6G1T9DyROkN6p4bzTVVs0NFBhdTImw3nIQGr4neDvp0x7g7nMZ
mjWdTO6D0yq9kSAfofWpD1paVr9pjI/AAiEPiwfvS9UJdYVLPzujbJkDadhuuqi7FpYFrPAmvPCO
TSDMwGZ4JVKvwaflTozQROb+CwZLJHKrXmj43er/vMLF94iBaTTtZonP6c9/NCla2Lk/s4Y676JA
wYzeSw5TO5qD9xOZIWh7KZmLNbNK3RBi7daAiG6qo05BLTGbbVtqch67flp7afwLAI9ND4QqHZyG
OHqdH0ELNqMUQX/Q73EtSIiNGwPFRUnfjdxHt8Nc+T8vfWKUs7xQU70lVSw52MFkzmqFUnO4pa6x
IseIHExlfLbT1ISS7jkCfgBfoKmuch63fgWDvRDOnSE7srlKMqnN1ZDmq7f8fpP7Y305GOlsA8aW
O6Zo6k1p1X0MMqVHSSd+Ne2k3Hg2dzXvGHnUZd2A/EJUUpcVEz25eHATk/75M7PP92axNhjJMzCY
9sx+Q60Q3iwq8eUbp/lxcCUb2cZ01xqLzrl1Y51Ga+iqO8uUComst/WBAvoWuoAUupGD/vNQJceg
GoxvxP/Fn2HrPzCkctpVv2CQfoosKYe8VfRuehTPO88gmHitoZ79UDkzsVS8rF8WJKvoQCkQ6wER
OljsXQbCphcx8t4Vg7yxLu5YOpVlNDmhgeNEs63ei/4idiNtR3WM6SsJ0ddxQvaY5+8OaUukDE6e
CZVj7SbXHJ/ofCLfnu5vp0azR/h5iQQx9q6z43hGg25WFiLab8E+b6O+C9LrTOZORH1er4cSIItx
sWJiDIHZZnqn7MdZ5ZWBTwftjpbLHO4jRLMcaFj0rg62UrcUJmnrqnTFARUPjqDJ6FkUrlGOlDH9
UvAL7KXo4gaAX8Xm6elGG4qRqukLWfgppkXv0fpWjeMV33Dg2FzBM/ydx95C8HWTvocBI80ds80x
RlZD1lJxOSJuBvTVgg+8StXnroy/fWCcoNQIQeQ9DzZdSQhdDpBy7ta92NvOdFQVXHVB6Y2mYZCY
dRvOCKJWL8VcMh583afoAqHqcL16/rgLGjkFcLD3th5yiEioNEMP7La0GDAMcALbXEDEncMkSNlw
JsXcu7WB+KrjP8PGB6ZgptRH/f/OY0UdTA64YtbKZev9PjH3wMS732wFwA6KgSLm/4EPUWXMVBM+
0120lgx94ZtPhOKMNfr/ejmG4jYmIaPSra1b2zdJRM8GCra3l0ZRHf6ybTro+OYYOkrsV5p+DwgI
BZxvKRsWwGSJ9p7n4qSk0J7jUt10jidsOr6c5K+RWGm3lRvxD5VBLqNtsxrMtqz8y2f29G/0AD75
y1twVGiFeJj0JLcfoh1oUhvbLLJAz1JJv4iQvuNLOAuD1gQY4ihNNjjg0t7GYAYmwMDa4clf1msf
qykXg95SF5twDmoFD9qSzL03HbyXrdERvylkuyUkgQBOAVFlkJFvSYJ6D8kFpr6IubYHvvyIVwhT
lVop9eYdf11UrW3psPKVy8p6QKzTpVqz7D6+S/ZS5DU1j2x5lkijNHEhN/6LfO/vY9053f8tTsSB
LOYMwKHrAos1rVoycyeAooJRJVcoHEPAf9MHEZHNWm8NIE7Ha+0pyJlVZcW7zzGDbeSyJXpJ3lIO
qJe334QM8cin064E99gufTx8ReZYn9mrXu50GnUF2ltC/3T9khjxdYGlmmJw8kEIXYUimklxpfwC
OWrvWMiUzE1mT9trlPJsxoMy2Alk18FefPM0buNlazGznrCDe8BVXczsAJsIvV1fk1ackH3igJFy
pnRR7DDzvrfq4hQDjDha6M4skWodPHbtDuwaTLLXppNTXM1DgVl2SqAi3DFL2I+LeArw3c6KFC9x
jusbdASJyuR5sn/RicSI+AVG0NvrCNqhqu68d1pq+eGfW5LlwsMTNJ5IaGDHf2IMlOZKDWxr9bkQ
JQZNCSJHJhDeiVuXXMH1yX+BCSHMTCePYNdIFK0tYX+PFXBky4GLKqtPkRA7EskVDh8kEDEQAQtb
R7vXILotgeX8TnoyUoToR/bdhbKk5BHV3C9hM/5OfaNUex14aXEUc6dn80AW9TbhR6WFwo6PkbXP
OCFU/wbiuAbaPCJWnEvCztVSLufMGl3QfztwVgsgCy2TPOoU2LstCjCw4aA34q3329b8lTHBiWGT
beErEFs1lj70DhsPTDGI91hmnM6Gf4HAXJ+nm+hmsw2JiEuXnvJWtrfO8ekz4da8hH5YNxWZVzgi
k4ZLTLQil7ZAT0EY4zjgBefe20Lu7ZAmuwXmlwrsnDnx3LhMIeXgacrz4eUVbsWbxsiB9Vb1oRK5
PJhzKrYDcCgps/pZ2JNMwlewzVO7233m2wdV87MO2yZmeWgc6AWhDWRfQY05gO9noN7aiInqZB7V
MVJxd7pSLvmL4ojJJAZPq2yBjj6X6nZaGuOf4g3kmyVxIgnx+cOaaab1NGj6leArRCRmaCQVKmqB
R9yZjBxWPxZgeiEsb4qW3FTBp/0c6cYaijwIgXz6NmmWfot/n4yj+U3ZICEePO077q/DJUjtkoBz
mfFJMmr7JQBr69kKuvlPzGjoQHgZcVvOZ3Vs4gRa8DleaooZ8WlJqfvAGgxMb0VupKawZJvDSXc7
kwqZ602GLeMHimKGKzdWi8EfqusjcbcB5S3YkBfZR0a5jhwnbMFV1J3zR1+MDolSSadU7ha1Ew26
GnB8wXFoh6AIgjQCcuG5CqhS4IMLQyj1X9fa3kiE4eWY5mlMfdC7oQQjSNwkNoRdWpYrUfBmGDLL
JKVhAsz/ZzAD+sXjMixqsaKQ2VW/fpAkdPfoF74IDU02irUOTfItOzjL+Dy1vNYaH617QE9G5ttk
YLQbZz0KWdGXUc7CcBvu/KEtkTR/q8XdGLETq6BkP4qI4GDoo1UXubPsOOmhX7OS8CHbKHbdQFNe
uZQpgp9wrrPlJTiNLZ3UiW4jgRaII2WU4KreVPqpHmPieiwYP9BTrDvENAQqoLdbqxfoutcx4rGK
ET87bngyiPKncu4hHRNlooS/NifPIt+L6BhiKkjjltJ9wRbMQePaYbHXL+iBKvVPgar+pGRoW4xs
zRVGKbCZ8AGuaBi1OdLLD/QKa7y4hx9+MtRtJ0Tj8v4lA9L0ioQUBZy8BOj2Q2W9q954y+P1ZA7b
7bKQQvoezKR+B01YuHsp4XcHvmfCESwj+w2yZOnkZ2/xIIoQusIqRMH8yZaZA1R0MwMrfwjfzQ/1
a3RUNkUuRevZ8YPGcLisaM5k9BcWsc6kq7zKi88mAHjJ5IMba3EAwdPWLoC5YIlNCE7ypdhHN4uo
lZ+NRIF7UGClf73crbBGaw4d2OY0q9CV1p05aS+NsOQcwh2iSBoFKLRaW5bpwaY3RPq3+j4jdKon
+904Kz63JrqaIdg1KVnx+BieIjQb95i7t/eLbZwB31+eBlCkx4MfGXK0PqET5iKS8rubwxok848q
bo9osE4jRYcjvTjpvbSJYH/l0vBLQ/WVVaaZ6LadAmXOQA60+PO7jnLycVNBcL0GeokHK9jB4q6k
SvtG0AsMDo9maoBRR9h5IAD/x6pnT3VLajUOM3nxqLwRn6IUSCBrnC+LIKs/2B1mTTk8owGVfv9E
y6mEfIE/6ZRaY+FcP0TXjEsmFh+9P7P5RPqflhqgthz512auYHaxS2QRYCINx8hPqHVHgFttZDpp
Dmp7OTeghO/S3uMHBKtjo0Fq6bioQJNRgXY6Jb4lbGfjeGfpMm/IWrIRT0msGoBlPVN64McABPuD
sRmZgddZc1KPt3vnjswSolniJXJepWxKwTilTN4WoEbGheoeKt2qSBaaWFtEf/Ij4NjyowHamL6C
Td2eonMZmeIDLUC1eswtbAZl+WJrWTwzXH6CJEBxNVHK2jho7fNrOoQbRYII5o46d6ha1mxMofAi
bnYhZt5Dk+B++yCni9tn/j0NV99NO+Ofva+8RQSHYIDTP5yd1B073Yx2TYCcDzsMQ0apTBoe9T4j
xHKksVyngU21CZoFbUPY/rODR5noEys0Pd+YYfwGYamUfZDO2hHS7mIbiyqyMCovVfJ5IF/0Bqya
EjrtL3l6k9Dh0bShOzT3sAX6lqm7M6SOgIn/jt127vTXdLDG2ohqYH7MSbqHrpRaqttf1S7ufhqD
3MARj5W8D7p+SDImwcC9Xgu9FbQ/jEYwGdgTj2A5AsrFr4OrzRkBsm2MNeRiNGmFtQy63bkLsGOV
hNgh+dgR6LJ75y/FQlkEXOEViVmJfmF/J8IkLgP6T5+rBU+5HHK5riPgX1Y6Ud3nJjXq6xrXalc0
wvN0s9Wkl7iDRFIzdJ/737afdp1tYU9DRiGNO+1rgK9Y+DA+IeX24N8ozlqRLbB/c+bZVSMSpriE
iCzFsuLiAfFKTiBpL5Fotia1hY/eupNjk6TjRHPvbBPbDjjaesZuC07bdWir8G/7WJYLDQE+yGDF
HYiKDJoizgJCFS/4AQAsSqWeVP4GIOwtyOwe2lp8zcTbpMGXTg8YB57LPjO7MFgryvFNjcbeRquN
IWWPU9FrdZqLuHaJVW9FKTz0iuWp59WWjKTErlhwUp0Mg08lISKxCCyPZtsvQqbbqD6A8xsv8mg5
ZDIfLd6bKG/PoHZ7cIeQD3x5DMc/uT8pdF65HJBDdoWwUVQemV6HS4nQqqP9Wj8dOSjIlpMkcDvM
onOCom46b2xyfSIY+ihfhliwMZV5J5z4zIV4m8YoL1oVEdRMGd9Dwlr9Rtz4fYDUiGAKo2HDdz6U
ZgwSBpUg9kmAkaGV7GsXVH2eFyHhmKX3YGrdzVGNs2YVmYoXt9nF6+u4kIj/wZEHQctlEzahz+Ni
mRX2Xd+kBBf3tu6WLGyRMALWKcm10kDszE9PTXkWoxW64crCLatDSSM+SqRNzLGS+I59F6wjEmCZ
8m+8mRCBeZbcyzPvSZn7n+Fa3toO5C8sOEhdjbpV7A+cZXl7mD039n6HbLX7uDeKtSPoWYEn/PQ1
bjC7I5PLit0o+RDME01BXRMXDilGDWZ2dHulAXmLk9dwkiCDjFvC2YyQdqG2i5A2as7xJYf9SGKN
iJ2/6dt5O0t6/C9v7M38U4jklXBoOmhCqJIHzBPMYEQROXPgIKnEKc9ESguW0rT9NtMXPbJ8BAOl
CNHmDf5n4fwrLctlIujrISjmxf8GJJVJyJ38pTd8ggbq/u6EvmhFwkKUzbtV+hwcDlXuXs/1+VwR
RyGG/2Ga8eW/mk9fh7eh5bw+O14DR+Lbxmvb+CdCxV6+xWpPxGJbdFzd/zVfg2GpneMGQl/ryUPI
iFFAyb48hOzrEf6BMj+jtr5zdO5oTOnEa0L2MqvL3to3G9BZtr38v8wPB/g+wMHfR5pfsDIkbsZ+
WmdoKiWTv3Gu3KmRdv0bu+8sf9k7JS1SJ3px0btlo6bzAfqVCvJi5ADd+3mFobJa3Qqa0V6SCEFz
62cLPaLjm6Lbm2n61+c6HGI9UqnlFavN19PmCiFoYlgNRmE/qRxfQfPOkHrSUS1WjpIvrpA3zLC2
NH8KfN76idh8h3BM+Ub6Il+K0RsfItfSXuQFCF2ddB/t26ihMTh0RMyuPUdzByE5Gli2UXJQjs7h
pah9/ZhsjNadO5F/BhRWJOp98z4EpOO+CpN5pHjPHTEMyXsWoMVaZOkbbncnIs2782KAZtVx+azK
XgBjOz3hUrzMTlEEY3q5M1lULU45Z37Ep0XjUz1XGJ4P5D07Xm0RwmRr1nK1FVzRW1YKp4KVePNm
dA/fL8SlnU1enpU0AQx+5I8wbf6KEvgTCW6LCDxXhp1esfbVnPsxXuRPhlUgr5+OKmyFpAsun5p0
CAD4wu20CTWvCUQ0nfMYY1vPKUlPjORR9Qzu48sDWktVLbYG6aazVTtTT1R9Lw51IzgripnsYUIc
86w63Pz5yb4fQqfNJ0NIV/zrZnYtNW5pP4R9zcb1lMvJ+0F0KeqgEt4lxpHKsNVGIxft+aXK9gaN
ZV0byoAf+RCWRUBoG1rFStO+Bgn2c3BEoobsInaGEs93O32Y212oZIqWJumhmrE496jBFMSo1NIY
NwbdRZ2tPJ303jLourAuF9g9Q/zCgCeGLbvhVA+xSHiIpCPnIKTkobWTtWP/0jOIujKn/FTCC9MD
Ry4M5282PSX4Vsnao+RO6/4jDoc4aigoPyg4JYkVDHga3+NMMhfP+B10r/1U0u/oegtYLIBMRuVp
JWsAg55HERJGZ7VnBr3whc8qFDe6UnZUJyvp/3C73ZYgdBCrCIdfGUt7t0g1TQ0JDs8sy84vVLfG
HO/Dovwa64vGbm9TeZZnUIuy3a1M5GpUv4fhdk/7CIVFH86THoRiG1vCb6ayL6DqcyfXwLJV2iWD
Rc9D21ZhhpC0N8o0ra7RakjX5T+CK9aL1O3xA5V81Tfh8tJ0G6ljMq7CA0Wv0L44wBjvCKoYIFEF
Pz4ycvZQOVGHDWlRjC6q1bz2yTSp04kTQIQFGJsqDe9p1nvuJ0zoCLtZotLFmt9oAbI4WPPpj3bE
UvCh1um4k7BOo4x2xeQb0BNQn10FsHfv/jQbUF7HrqZHXiXL68epsrgSgmGwv6zvAYcFGVgjio3l
EeZKj/aXIDzusaY2XqkHIS+4y8g6tPv9GBIUi5X9qDz6nf9VyhRHslG6OzvDhGmTnjYKbQaTHB4Q
5/905WMuY8dTMzP+ApV3Q4YfyGyVBAGauc6O4zi93obIZzF0q22s+3WMvuqwy07hEOXRruPR9HJ9
e7FyjAjW77k7bIMxu1SEwXsKluePUnUNvHncRQHj3bPOgWy5ekroyCZGsSfhTE/iKelncTg97bPs
kE3Xr9tEnAC5Bkd5KnNCIKmTHEluKXSOI8Ocyv1+k6LTrNpZ2znHazn+RJKnoyllpdCVXzlsuEvF
1DXNNO33GmYsLeGgpdpftgA11Cnln4+p2ifvf15hq8Q89DlMhRD9nZT5ECgOWXIus2/CuIEXnygV
vwKdF1lqi+IAvVUlM+2NNBWME4RXmYQYKqOqQ3no0WMF6Sii3y1XyQgm1nKwDqKhQThTkSzB1u5v
A5lKVvbf5B4ZL+dTLTqVhgDvLiPFn4pm/izPrZEYvlhT9D3+PDRfTFasv9DRzAxi3aiwCVt440OY
jHVh1cnAO/sGKIHzfN1bh0Afa16y0a7m01LWPyumaHeWNq027pW3AEmoFKK79khP5FB9h9M2RRik
+Zu9ASeWQefnwzGwXNDPGmHsF+K7+YF82gPfmMEjtkZCo0ZU2+p2+u0JTeuj6iS8+fv3LMciFV7O
ZFSuqcSZP3o5n8L6+jkeKklfEJb9ud0NX6u3Obm4rYv9nBTQysVFz+G/a7b81alPLmYun5sulL89
IATKSrG6SXQuPuBe9aOgglx8Wn+LySFKc/v7i6Sg+ajydp8iUaG4Ok9TLLSM/f7DbZWVaYt2MNgv
F7vszzKVxD4HhO6zbtrDfA7dSf/fsseV+/1mWpuZedBML0sON8GXGvBfP5dfPZLtLS3DBlI55Tpq
DQl/aJxfjUY5G0Qbmnk1JN15HS7idJsGhlwAvGvy1fxHh1dt1YJ+NQeLdyXbB+5ZdDNkXdaOd5Zp
OMGvKz23ms9t25Q9ET+u76qV/11DdjbShlVtLWVMwR9a33R+h3nxIPL1EoM6dkmGjsgUVlzRJEVH
vFTG+y4ZcS92nlSvj7ZXdGstI+W165paYGMXOh7OlUxgXQdmV99+tdoFG55ElZ2UNK8QlWIQT6S9
FmBvMJbI5P2VqsSNaABuMTzIcsTy0tfc24y2R7xCc1uzp3IVOFpH1tKduLRxPOkX6I0vnK55YCCq
m3Z7PMCmtkT+dQlhZwJGtWBCeZVdW+fK+XaxQOJrd5IlssL14BdRKIW2Ld0dTjaFL4jdj6t/qO6q
RGHJVK7ZFaHxVntXK5btiIZzleV6Yb7uPiP+iknHeIatCVx/Ga/+sMM5tkmveceZ8E/E1d9y8eZV
F68tr6Jgg6cs2bOBym6yq2HzmxW77I7/bWFd8LGYm6Kwn6Pe+YzSbMTDSODu7wQfwN01sJAeMV2L
bwJB6LpU7aLyiwzHszEu64PleskT/I1r4od+jJry78T/3ykSUw/M1O4s+AiQ7zyanbRwBAjgcHpo
J+iA4N1PQiqYkzggTnz/8JtQg4gjPT55zkFUKx/fENyNMrtVBpJCMfn1ov7w9DvSqytYTCww/+Su
0JTTvruGePu0oAnmX5utVMKpal6GkkWQfZHYI/5g3+hr1A37FefRA1xc7mlyUK95J3rdfo/Ag4s1
F/ENVb8hrDWxutp6Myh8kaS0gg2RO3oy1GM+JqgDk4Uwe9RqslVE2ySyhvRmchFOUxj0H9SSyaZf
96wgeNQa9GXGdv2V5wuTmvt5/oH36Hx4JXm0RDiV3QkR/BHt9sHLf2t5uPlWg1mBy+OWO0E26ygL
T/vpjNQPHz+BSFqJ/uNobFWYHoSXAHEkpbNxE1m3HDjBh52cZgh+E0aqy+w47FB1YjZPxIvNrW0m
ZixBrm2MyvMklUsM2xdgF/P9M5xR++boLki39kr9se5EY/7itKLiMHaot3ZQXRnPKYQwCkOgRzJ9
ev4P9Ali/UUwJ7wYAs3ORy/eZYsBgV7ZqPTurtYIN0trXS2uJTkM5jPIPUpwq/nKk1RuGxE6qOgP
4Fo1Z8bZM03FgPQng+3uqIF0ATMPx7lfjTMDhuTYKMDhM7HUJT9WOLvLmiobyCls/MhXTe66A+G6
I0Qhu+kS8ECmjX0as9+61txoARc8EiIP4Cp0++sT/Xc4Gx5Vk1FhLetPAlHsZRfQ3LvDSqlk+4JR
Lc286cW7w7T2Q0N6NIT4jNGDySosGmVtB2xPZRTGid7UrZsObpNlwmuw00BuVK1eaCCTezZlWlZ6
eo9aabdQngGM6tdLLlV0pE5XI2UvxIZj6AxxTxc5Bsf29UthTvXp2SWy999H23mHbmaqQcL/AM6b
fib7T2MmwBGcNbk+wn4DNbeOjQtiazgsqiMS+7I1cZCd5Vb61QHQpSJ+6htIslgTQKS45Qkj8cKb
rkWNgWD/scVtjh4D9i0Pmfis9A0YDw7xHsk/2s7UAqeM1u87+BdS5mYbS8yU4E+0Me9edJwLF7h3
75XbdeH2hawBDcllVqrPqE7HEZTq9vFmRBrRYJQnQICUXrVPxehbcx7CoJffH9jJiXvwV1Y1MaDT
F6wlyswvXN6Ha+wpjh11rLbgM4avUFdBgp+il4d9SPQZ8JrDNlv9mIN6ONMClJaAKgeS5NruIgtb
bQYY/HnTmERUQpyRJBff550jh/6cDTl2gVyujMm8IXFLq4EtWOcCY9K7GWtBtbd1WMRWJWXf26oQ
QJ42eX0qYcqlNtgsoJFimoBQ1psIlluXkAHk193X4O0YmmxAsu76Q9EA1DNU+bX7/YQynG+hzWHU
Tg3vvPRCSWT2AO6fUGDQc9OQGrF+YEjDajeDy0Khxby9LEL5ewSx38Yuo7B2FrcgHl+v+SWLgyPt
S4CorAMrIPrt51ItfMcKSZmaE1xcuURIuet+gpY2y27UYaK5nZPFMC0q8eFWIpL8/gAdPPB96O06
WbW5DAwjAs9cKCcFahYfGaWVzimkhIAy0IAx6C+aFcAly+BjUTJuFPZcgtVMuDX331efwOaEGyyQ
UkrZaTxZ2Mv/t2wXRYKMrgtSB1U6WPHDHgdmKLACEPXAldCgrhMjCkwY62rU1Eiox1lVriiHcTf9
TdfJ0zsI180EzjytZHlx+jjlLQOltxR3i5bQPoiRovZmkxilk91OTEVhjyMFBvyXW56moRLgRz9Z
dEpi8ii75vj7mo5Ubn80xcdOHDxSh2t9Q9fjIVySokiCtTHgi1kV1jiyJM9O8tefRSlV6/VKj2eP
pNguJGZL76okZkCWUVx3pFisOYAYmTpJMQFfX5z4d591l8zvsXjj68h9cyq/iuvzzmLghDqu1vev
Q715Uc2/OBzaIVnxKez5HZNkqSHnTtmlL9AdbMHE0Zj72FEUy374pXGkBN8xasOMsAaK9Kb6MOaK
fDXXUWUIGuxWylFEG58WmDfQxsWDkPmho4BVkiSwev8ypAMnzZ2KYfDhbd2tloUkV9Z+VimGLZHL
BvC5UC+dYGkpykgyq5SAv8Fp9WTPrT8s/SDLLEhS49O5hEHj88nBW/8ced53WfXN/MA8gDTZlbYT
a3fbhyUeOD/tdup4tjqtch+FspSR3kvuplvxUH5mTC3Dd6d8nHsgP08uQk/qzaPgXKXtd9ESKPKl
3CcY0C9z4uC4BOAEJLMKHp2datqM8g/leQapKpsFHhszFdkG4Ad0hyN1TT92EeB31rDRx9e1Msya
35TINJyHH2fnloR/LOJl+ol+34EhhhtV3pvC4KQqy4RmsBUtlE1/l6tdFse5P6TN8g4add3yh+Bm
DxWNpajZ6X+6s+RBbNe8mb8mJdC3M2QgSFCKLlkvg3dX/x+P8zLtIlaKO283QOKdJrErFPbcq3rA
N+PpGi2yEHSDtxtXPpUErM2exGlTt4wGb40l58rvWAG+P4vtdA79jsOw9RQlNaVnAiZHbX9CFGbK
nlrSqiIxGk/98SgbnKJ6+AeLMZWB83pOfb+ky26xXgADA0yu2DUALp3qVnAYfX9t727G103tDKwO
ZWEiUaqPXGXzq4wbOoKq/Nkx1Bp0/8k7wHM+Yq66sd+ZC5/O4e4HNhPV0flVeE24BnFP8Bc/LrnZ
NE/c/Ov5rZjie8Yakr8saErlrfpVtGm//+M2lC6zdiCYmV9QYJ3DwAxcldLIGmzk2cH5hnkVzKtR
hXaobsPOtnnUFbBKJKaa641w+iBuyPWqzMMiCNoOLxq9YBwFl4LVKDzVIM2nixSea/X16zB9h11O
XJgJv1+XdKp8Jyhi0HcDW2JxXocF4ebAZS4XRn/KlFTnZuz7MksaFl1WNuCgX1pCyHKc/w+xRH4o
KRjpTkDH4XKV6DEQjqZlfMsUawL8KTg/w/kfshsh+/vyfB6RCqZj+o/NP4BlIEhB8Jn9vMVKRfP+
MxsruVRqNJQIPKotfmyKdy7x4PI4xUf31/W+mJA4nlb4IHpZWO66B2cgt5ZCQTAYOWu6s+DyF64v
IzYpD52sIsdBEgQUBSMG8vhVN3D37feQf2lCcUKR5Hl7MAX73LC5EnteeRiUDvlI1jrMqMblodkn
+dbmSNj4sNj3Sm04VA5x9S+XFFn9zPBAN6sbczFkUgoIr+nIRKaV88MhNgWtQu+ie4cqi6n70arO
LNtTFeMJD6s1EWvmwfMV17S1dCrGMEXtCLK4mfF2VMlRZppAuLD1z3wX3sr1cQwgCY01Iuf9XZps
CWH43vSyrXTXpLql6JATM6YGPZJ9ks11HYWNJnIu+83lQx8mwGCTD1m5LIQakOEU+TbPEqrdkYue
e9gQBqweRL05xC+oi9W6WIwLR4rN1WzX3jP6F82Hb5DGBojbOla8ulVUzcRruDYlXZZZfqL1X9er
iFme5J5ORBkBRCeSdmYrONu5ItvP+Ne8fy7wyIIywnLiQXbDcku85NCtMPNPTOqEuj+ZhYywRSJ0
osOw8zIDkrWFz9+V//AfBjFKH9rAHUVNqFkgwalbaLwlUqPbUpqLTsbeXJkR/wgIxyUivaxnWbz0
D6Gy+LOqgdQ/0Eh0oSxwUW39HeC4J1bqmtRJbKWNyFdiOa6LMhuv7bx57UznvWu6QYr2RiG/fCb+
/NGuar5cU7DBP80hUCIMLqHHDx1oRZR6+I/2bv21CqyuY1JFztM5cyLkgirXxXZgQtCiNnKj+fQZ
vNG0zsOXQ/oxBdCRoPI9mk3hVOFmPfvTecq8JfIVA1Jjko83d0gbJF4YGjTLbf77UjkvlNETxifP
9CvcZ56cy5lsVOHPWVifvxIFahQM2cPHrWvLM07OOhgid98bRnLDbrlK81TbDJ1nOUUibsJ7gzfT
X/SMduqqyVt9H7u7TmR550KtSfD+an+ynuDhW3CEaPzteZ95TkQqU6t4O7FRQoeoH+02fA1zong6
bJLYd3dcvrLkdIejsCo0zt2XUOjmjwVJzZ6Zk6ihdzt55B9U+AZ3erAF+CPg8/tAU9zhHXH7ojuZ
8360rmDsHxN0OxffnRH/OLAA543BBKuYZF7vuBaVis8jzuKs0EmzoUEV5p/AlHBwIDUmdNJJKW9Z
6KnIJQDtrqgCxW8KYkMYCabw3YBzo7kAmvTXngrlF1j0eG4mSKFnysjZT0V7a0ixH7Cx6upCFHXr
eYrYiE3HN/HenWKJQ8KQyLr114QeKxq+ErTe7lfL1AW+hHPnlWZGpJbd7NksR0h9jqhube1FpJzq
TVf8UMsgPeKUWh2PviLorJ7mKaKl5HEFhmbETd9nohBdQB+B8rXF5hOanKTPurOiNoCfl72KVKJQ
oVd1FElENnAgYNVlx8v+cz3c31JBfHb9tWAnIgoL4/71ilZvTQLtDJOHTQAOmhD+lCLGf+B+VLvh
OGg9yviB/e3w0cbc/3rZ8gbRWPptR4A+Xs+uUJ3F5BZLM3XsC2P0+AF0Ox6BpW8i63o2xzPihJDV
l15kwz+3F22rxuqO2oyxSEzqGQ1s//5uALT8YhEYiUskjY6Cd7anQNnp8fYwQxmwaCWuclsaq4tm
pNq5k/UiwH7mbobo4IyRjYZkWBwzzEf0InGYaUG+aitU3l0QdZvs0T4YhSsYNPUwpR3gp8lwko6M
sM00exb5g78xFsKuwkC7+tbHpefRb4/3jvutExXPIDGx8kpO5wHvuLRTwDQJN6NmkYTkP4Z77WeM
EjQNuewIyy/x5aNAoaA9zJleUg13k+0SiUlfhO9awL6rXi1Rr3rIGf+xLw24sbgPsh2gY/bGoPLI
yNtRIjjEXWNCpk78MwzAwVrQJdtdS+2+bj2WTGIcnmnZlkpM8Mf6ap/TfuSOa4QHChexIIpjBT0Y
EmvGXyIWcZ3y0j3SSUqST9DX45NxVqZwsBxpWvEqemNPUolkKK8sHm8bCUiRpKlhL2AtGudiTOuw
rzyKx1F7bh1PbPmdOE1H/x2F50BtMKznuRcYHDnNRyVeyNzwjuM751WpHvO1dsuF9R0ILuAp2Xm9
Mi1Imda7oqGTW9PtpEwb6vFvOAhpkDxEe/W8dt41hqTaNg9QI756Ygf5DpIpPMzDclptEF2UG3Yv
EaEtz3Z69wiEplBjF7hlUqE6ulveLatDFcwc8j8gCXhZFV636wXEo6USVsbg742Wmzuk3iYUlhUR
sO0lkxlGxKGFwfkIbPKPa22cyg+X1yH6Yvey9OEOh+mPIfe0OOPH2oG8QJOChh6OOlya16x/OtGI
hPF91ILUyBTfFfbElQnWI1n0A+0XwBtvUojAcY3AN1wQaxLwVJuuIxfUgkNe8Ak58VcfHP3dwA12
Cp0+wjPS5wjPiCmU1rONcdXPzFav/o3d56nSoPVhBzrnzohgujBeKIJr9CoMHcPdgbyIectwXSw5
Q6GLMHmWZHfRxxfIzsLH4MR+oNjKwlWeenxhs7immU6OOhWivkpBJx6jv7Tfld1AJNYsvrmcYR1K
aBWsjQYB4KqNzi7ejeg27fTjNW+FEGc9ySAPtUd457pMcf8L2ikOSFf7iYaNTYo+Krpjpgjuv6+N
/m1x2DId86iBx0bzq/KbjmU57J2kGQKELr9hfRGCson4pqz382/8smXOWNKTCdKTffZ5up6+XHiK
DxzhcQOgEVqmQ6WFcJXm08g7iTIYAB8EKdXz6uIp2FKzwL11ZZEQXt8YoMSyVpYP0JzkSy7Z+02r
0zVKOmxKz49eAb7BMaDOJG+ZyVLAyQrhtxkWTV4D07fyKU/X5zD82z3azD+nbN146Qe6GzNQ5dGo
e5nP9eH4eKoAqEW/kAlDGXUd3zzxk7kn9PH+q3RKrweof9rUW5xoQyVptfExogX4uG5xKoLSOTxb
6GreDxj4Kpwr5BKCAemg5nxnlh8hDSuLIcL56KbQ2gaTgswtb086WvM/f942pTQ40Re1U0nyuwl6
Gy/cC2jicw4YH2KvMyvpR28k1oEkPM5ZmGGmx7ra/qd0MuIPTUJ9ZjoJl0NHjERiCXrWK+5I1K9q
1PRalNRxCKp0ljSXhPoioPgE3+MCNHZu3hEdIoBaBs8KgZJgoLdlKgtI/adOcyclAv0vGsQVHMQ4
xuTOpTavzyfF58r8ct1dIBkQez9xpGmObADPmFynHgpl+CouzJ4IXgRbuvnyIePbM/p7cLzG/FMH
vJWhIzh4vsC5xWQC1U3yZ+orzlIPR9I9s6rrxeCIXGXJc+V2iAgheE6J6zJVp1jYrx4Q6XyiPJMU
+IxtWL07Oq2MB4y8wFlPgpHw2lDwZ4cUrr28Kc2PZJogu5Ibe9T07qNPyenMMR9VGrPQp8cRwF0f
n1rlsflkaSilHOJn0uYytEp39B6KmmVEBcx0MNlbIEVe+6fZ7auZzPIftGLaXYrY3+nS9r6AcyDe
G05eTScJE2ZdOEqtcRJlRPqv+GPsdxDNxNztGvVV7V1ttsKujc/EYf1S3vB13H3d2pQNmbCtoaKd
2vflMuPPk22E6R3l58Z8yTat0mfV5sgwWp0LChICkLqVwYhQyxbrV74qIo90alFI5x0lnqL97Xtl
pF6Wqi6/BLxoN96V/wQ53Wwfg7sMAHoOremyke2DTxv0XYlEfj1PAV3NZ8HHlQktoUqqHOcUvsCK
ybCObVgwMjDnBCYBf9kJf70ObIsy6X7yvYcJ3Icsdzu69dMv5ewZFOfCqSL0QNqifRH8ieeiP+M1
mjdNLyAzuT4boV2bhV4mvg4i6+g+V5Gss0+ugQE+Lrj77W+lnsnujbsCyXPeHGKbaQvoVP/NIq1o
51H21DMRWApCqM3Zl+W+Uo/W0yiuI6BnNs67OijZWm+6vawpXUX7+Aez2v8CsjT7DPVPXAqpXwK6
ncKO+PIH7GJ6GMAILdOb8v0U71A5ICe14HIT9qnREeHxze4BlATd3JwuabOhsiIsIxkvsbFUTBev
R4e26WA0hHffCdINN1Vb7owYVENuGc8aMQpHAOgc5eO5a4zpbtKpOdWqT5MeghsqxVDFk5M//DJ2
W9OPPXXX0rMU/6llvyCbQ5Fq07mVKs3k7lpR642C6yPL5AfAKohgtNLIluFBe/mRVyye3sUTGicC
ELT89eEvPAK0oqyuG8LvVO57O0HEJizveovdkwzP9B5ugvbtTHrLM2czRsNKdT/X4yxxvv+BrvQE
dvFSyK0KJlayPgm1kjnUvFu+E+SfeCvlJxRjQGSiFJonSVW4/yYI0BOW0StEwGfjpMoExS7odcOc
luJTMs6a7HhHne/G96wPHkb0XE+WY0QUqH7yRvJhMX5enykKmjYaXEHm4Q0501WUoYijJXevoRIl
pyklkdnoLQcUqHzJxPXTZfNFBuxYQhOKBQ+2/3dzF96UPx0MRT0ZzwRNb7N9z/JWUCRzkZRaLSz4
w6w8gSi80B+n0d5j0JAKDoyMbqUTr6Q6Q5FdhGL5DZFxom82mrBTyPhHDcntePmZoz9/aqD7WoF1
0Lw74y8HkzumIj7FOdUPksoj+cUlXFwZgv1Ov96L8V9EanMY5ZvIWWHDNV9Suj4GGdHrSbJ5xFPG
gcvGw3ElkDHZKC3U4gXDd69A2k6YzQQzSBS8eac44eLy6Hq6r/wP71VDhSSCGYTg4yzx5oGKw7os
B8EV7F1QDzYiasi1thQgARANXwijHbc/wotD99DfO3wl61LDs3YIDyNr/w7pnfj7fM4HW6Win4Ix
iO0HJBuLGuXwFtjbzHcUdTeAhZi/P3S4/d61W07VdJXIzX6Voh9vdEZQdBSp2QK18vh05Y0AEaHJ
nedN0C8RFc6EZFrfS8C/CUSlcn2UnF1m0iPBmWtI1HKZKSynytth0yFk/bGIwSris7tT5WtfUS77
b5b8u16I4YqE/n6T9n2TMwF5ZnwxzFB6MRtTC6hs04c0wi2vmpDuT6F000hxbPpEhIVMJpmrnD/b
4lqzSe8XZc+7aBFFemrNzgHZ1s/brfcEuSiIgbaVztAfOriuM6oc8kR2Tyi3nFu8SOgH147zPNsH
fhKzaY/rCx/NYUgbU5XKeYAkSJvZZMjv0obyeVhMaZD/UsZQp93rV8fpMyO5eUyKA2ui/uctRtCK
hrYLpnzt503lX/eJrb0DScIgk5ivkoHOglZrBcE+RvDwisgMlKzQWSD/XCdStlJ9I04HOTUazZD/
Nyqnm0M5huNpVBhlVfj7yytyFgLuORK4HZxX44MQ9xqgOulQQwbPYsUoZFLfJV+VF1DeCojX3O4Y
BXF5kajwaWb4e001+OEP8Qst/sihV2NC+CbRHnTngIdBB8NMEICbcymINqWCidmFqAs++s6kdVgO
oHJy/+sOVLoGK9mkG2ewgju9X9F6HaiozmArs8oapuzCucjGwC9Y/7W30hRdUigqfZc1QktE0KwS
WVDew39uurD/1WtrcPKwTrWdhpqt0utF2fmIO6LmJ/NFG5ZHLy+htNXcuGPcNcIlw4vU/A64Iw3F
/WkCOgpZRTkqd6YZ5i+dHepqIFfEx1W4zKCcSaOCgNrwC5WeOe+Kx24oqV8419sFD89c5spWGUoY
8EbuyS1iJQIqdDqgd/VB2uHGbgH3cK81MGiIKcDxmLBsd4MLQDp6Mad76pt7OFfGXt4VN5aYKWQc
m0c/hnZQYZ8A8NsSoh7qHk/Q1sssYwsl3bMLqPLtCAx8Iaw4/ioSH7HbNBiBe9BgdRZnBw59WM98
oRfgjbtV1eGEnvwraPBncJxFTPFqwtmxaW1GIuiqfpWtW/a04BtP1RZxHbGY3bZUF1ge+jv2dZW2
qkirj4xwx9EyOhaZSsSqi4uJKgWPQFH6AlZ0iXrWddmuKOusO3MT6yJ06PKFQdlFWRrEd1qVz35f
N8UP96SVqy9Bca6pBxIDdo3Qpl1kPzvVllRP9Dc0dGgzDir2sSxnQ7cMC9Y31jSij5dZOl23Nlkw
johoVJuZYx3os9xRulTY25cD0E+teJ9A8GzB5s7MZ8y8P53BSIGsJOObtczcorxwKb+lqYojkRB2
XM3wNJ48TLqRa3/rK87aN6MO9qcKNsiRa4ToNbb0zVrZvota8aM0+OW8Dcvdcx8iDuijaapRM62E
+fRQ2nfn92keXVHReSEaQKr9rwBZmkP2UoYcpwY016s+N+MEbjK57okmNghPbY2h6Jh+6qV409rn
2epa77vBmMP+qW1D7Tp8FLwfhdJGxItqOXb74qJwxbxjma+0fWKfVKLLaHQZGN7El9LE1YRlosHI
1z8UfD7fTGwX7dybiPwiIrUyy6HjYU5TKPjrw7OIZGamenMxm3mC6jElywfoSil7TGrzDeDOvFLa
ttXvKhAiVQRZtHar6Riipnzm1s+BlWCjMKH6FYcmpb3Wqebb76YeIaGDmg1AROeTjYT3xB+ZJ0J/
+v01C6lXIbzrwV7sX0Bp9kgB+qM3bIrXxv8Vv83iApNabrFe+P6k2qaiNsmfHEAXiEWmfh6JqN4T
qhYB0qf+rDe/JwZcD4Ke0vzyiTmY9chATiLKzkexqc7F4tj04ifnwMtnTze8n81OuplxKPPHoVbX
Wm6bsB3y6yYSgcyxd73OUNQeEmegZBJpB2vUTsQBesnL2b1GCFZXushUPV3fkxGsjhaEJ9YdNC6n
g0o8SPJjA+Zm7uGzL7WtabE/Ht7Oomziadm1stDBtoyT/KvwsgJncRr8bkB/MNynZsZBX7uRXT85
IAoMY4BkK72sixFomq+WIyzcLrUraO4C9/oXDBMNePC+TiKKQOj3mAjvHMkGpzp/2bat3yekA05P
9rzaPJcjl0DQ3/WePYooqlI4Oz71wdJTJVu75Hi9sMDr4Y0uK00BjretjRbSzV/nxdlXZsJpLJMd
ihyoua7fagio8s1amm4vysP677H2Ba/BmZjFP9ity5UinxaSAvzZk6hKX+1fUzMhu8UYrTQW9FjM
axx7lzMW1mbpisOZ7O313pt6Gvc8ujCLvsxQ0F9zPOethXlXZsOEehZSR81UnHNKJXQTd6c7nioU
lQ0zvuxvFtjR3PgjAwZsda9FS7FGUoAsbryYeqaRbnioIdptbbtwsxXy4bgiLAJqujZDNIJ9kAhI
vWiqlt+9er0OE2d/tnNqiHXoplHUlnZ2Fjgt7ls7glNt7Iy0DMnaQq4RY5Qpja7VAK3FUf0UwWAP
5vtv+OFVQf8F0RlaWpNtkqSrl1okCnIsNdS98UoLCWz5E8JA9R/xzIkzw+zeVkZ/9SN6Pw9PDQAg
rRTsB3jBktT9clFdsU5Dx8Xgg9eit0pkt7PngT8l6pXCQJvqGKFKS5gewqvG2GVumwfj7YtmoE/k
hlTu5HpS5yei+D64bMmbVzYww3zAVNr1yLv8Dz3/TcFhQsUIEUyIKxvPLJ0943rQJ2/fdltI577L
EWstXeBDt5ZlcpKQOFQn7ZwB9cnZtE/HcIyoobAM7wCH3WTcVml/pe18OhVcWpAoa0e7VF+SuLXt
20voO2UMfaPWv3RF5i6x3wAtQJ0+m6e4elEoW8ciCNkMwvmAc/ZHGCql763MJdDl3/jhMI3HBRDa
Q65gnU7UoMEFBXv2NArHfVYFkqrPvmru3X+l1mZIy5raVegmeeeXD/Ov+Ur2sBH+cjFs3sFjd2Sl
7zJY4dDlYQK+oCth2wEGc1XCXeDOGY/pq/AZ+i1NfiAY8grUw/eYQVSRm0usttE3/lyOOGf8XBqp
/0G3i13sJhLsBoA7HW0iUzPnQz3Y4QGxKgAp8AA3sA7lgNVBLYlidEXvIms7fHgr7CHSsCNn7FU+
r5NDJWhfT7k732ffM8OIiNR3sCoWOPSDOZe5kkj3v3Gsr6qTVdq6OUj0bIHDTF3jehHeIOnvqLyC
RuU9ypCNrj0NUP3Pq4zl6iNplNrHt7sf2PPNprB/0N7Gzq9UHfy3K7IHmcKcrfLK0KY3t9qYOcYX
Xz61A5SLoj3cO/ECZE9IssxzrOD6fEuCKWjY8fFYjQi0iNvUpaWBCO+cPYgQGuSUGkMB0+vWgYSj
jDYssd3Iu9HXAAOR/K6T4Kz+DuYi2qjJ8uBSZSJhHwGvOfcgRDYzh0QKe8Lnq1mPfc+H9t5fH1Jb
syzgW4+cTAv3n5NVMnoBsLV+wCfVpbvmSiPz1fsHsuF+DtNgXeLE3WGmkIUZ5wV+IS6LDFH1VVch
8jmxnB8RSKZyY68qYB8bDm+qh/fuXtYGXJMx2gakjntNIw90OigtMMpuBT12KBKrMOpI3d+x1CDx
XKwfeZ51BF7z9saSgPc29jvef13vsNAE7O/qIPyE/PY8hgK9CEvhILMvgTfDYIkxiqoyEPbbfaOK
JWL9eKAl/WDjZo3nJMHNVHMolm/HBYbNl4LJsX+l4Tq7VwH7eJ+pVx20ftgV0kIMlZpxZZ0310r8
BN3CuGhWVX+2d/wqj4r/NKmYxWVubG/xw0YVkvQIt8HDbnivWuEpo23+KyG4XOPyBYy+Z/rspMex
mnNkvzIGEX2avDjGibBvGdbGG4Hd73pZIn/cJc2MLPxdF3tywX6/N5QQlvxAogVEndNVYZrP3lhT
MWJUcMyIYfe5xtDTGAhI0M5SdH7dW5zosqV9o+Oce5Xho1mRT6EUV239Cwk3K7MHifToEmk7YQCN
R4NtZ7jfeProz4lSOmQsc/h0rD4wqD++7eooKURAVn3NIifvhuxG2CAyAfnulsqXp59hXB8uyQfT
i+CB/boESBi+Cr/J4vM+yCfxHxGKdmTEALCcQnXYtRT//4CqcakZW3M2mliqKf9TtoHDLiZTq4VB
04gKIwVH66OhXa845ujA0X0T36y56H1rTkvUAPvFWWdy1jc102GXIGYFgq3JIv/lthJudwvLVbOQ
b/6qY83wKYEWVWN6OBSpdp52/cN9N1+e9TzSYIJotcuA/RmM/zyc1zlmhjPY6iNbVSPaIMNjcz5V
jUdcmKvTKmrgsJZQ6J4GPTHvQfojkZloRwoxBiV2v5IPE8WsmNCCzlD0ZSoyJucDxiWO6vW7OYIh
54CCVfJ3xAblP7s9iWw2Mj3RDgYKODo+43yqD0o+IeordC8zjipyUUZDNTFrrIn/XkAC3tnBAmk0
6aB4p6HqEJb3sb6ViXAUY8gp7pKpahjUm8CLvWX9P+F70HFnK970/YDXcy109JI+pTDVt+x+Me4z
WEGT94uCy3LCApGk0f6cQlF5UmIQBmrZY31qjJfdl/xhxea+O+leonVU9XKOdjBeXLQ/4Jr+ochR
eIM3tWnDb5eZjjsG8P0Eq9s7vKuJ7uK7/tGF6Ajg/6twDltKyoDhn1v2EI2AU7NJdbEd6bYdIzEy
MFgrW8G5zC6OfkfKK4dCssYS/MpjF07T4xcESfDOx+OYjO37MBk+Z2psB3GAHPmI1aU/JTSwPy35
2GqSe6nF1XMmEs+0J2Lua3Gr9GlRY+jbB5YPQaMlrqS2nZ6ngN/QbxBaoNB79/DZUAQp3z5MoyC8
LAMCBCgT1TORakj/3X6C1xI0pLOwp2dA+fEpKsjE6y/fIymg/7YuT+/81usglmOs6gsl5lpHtXER
GKfLCAYGI4xnMXv0eIOH5/yUIyt83xPWazMK1eyjfd02jh5s8sl9IiXr8KP87Xc0LJw+aHAL/P8I
yKveXYHghu+n16fxtv65doY0bFL8nCyhs2ltyjKKijrJrsPcrQJmK1CsuE24FmA0otsnyh7oEYUs
wrIsOjQqRZdEVknM8XzmB0PETFusgRZxdomOFX2R5LyJE5DKStlyJhNyElxd4OrHgn/6DxbMq5rU
wRm05rLVwFK64bZc76rWfG4hLpqAB1FrO4/LxXY0XkxvW7y52kJjMKuFMaN/UouGqlJSjYIzsp1L
NWxG8JNT5EhBLgChEPUhJrAANvH0k8s6wbBtg4YklyPLgPTV83I+GO2tGDGLe+UGjOH0cpARv30z
yPd0xuNmrZtGzszh2s1rJjGXqOX5JGESh+mxpzKvKH2GeLhkAAKBr8ubKbeFaCQ8QD/zkw7LSvpc
KwLB2v+zc2ogPupZFRmqpUuj1zndK+TIRr1QmyTh0gUwjPddlPBOxdiNcHQWVC1q6gBK3kO6ayrR
5+JASMzbJzyprDj9cb483yPS2RxEQil4ZvTN02byOr6QpIIGDJBgDvh8pYP3DvUFddytTCjQVey7
yQc0RurSJZ+okbgyhuX3Dz0WTubtd0SfopO7IA6u2TwxItyxBSMyPIHL9WTXcVKuk74Z2oxWdeIY
10Dfo3oAmReWoj04+by7ShH166uuFjKU5aE4r6FpjhNSt0oN/x0bitRXbICA6hisBA5OJ25Hsp64
T4drQpedq3hjMabOzs4Py9beh6yI7KfKCz1npIgjiFkN95uEr8nZZam30FJu498XXYjE9rXXwszt
Yb2iFpw7k+0aPRPTnidHCQ5TNyk0/QiKGKTgC4Q4MgT81MQjOej/zAgfzpN1CNjxEjsRsDOCCipI
WZtNAOWG1otIoUy/LrSzUjOyAeE7jBuW7bQoFiAVvZBTyw+tnEBWGHf55qMOVcf33OdtKFhkZuHw
JrR+/+u2tFDqGqYE2p28zTMpdH47QnCXgrF9wTcG6OqQzBLmfOdBqQRuemaDjwLQz+MvenSk9SR/
2hx9x+l5OM+ge/yM/GjlC2NZWq+szZEviwFXfBe3ce088TJ+sdGwn4RnHQ92OiMc8tD4dMqwDRMp
4BAA2WRHA0CljRXkl/xVQ2/acMShpMt6ZVnORetHGKrVFLFWtukE1WnBJru6xPLth+qyZo4BySYV
IGYyU7bBQIyJhoISMo94yfZmoc+gsg0S+mCZBBOKnOShPGZUdHdCv7iBhO1LYJpSgZvJpEhOm5Gx
wmWl2FcgiTI6wHe1pdnwPEsWishN0mkuzatgI+6Z45fW+WVSw4wx01cdH5X/VrJzEMNHDR3gT+kL
D0cMWSc7nukbicP5lIfLRLvDG1AY+0DjlKfg/rEQPQ7/9MI2Gf/6IjAzEmHI1PXZluXouHIw9+r1
LMwbyc+M3pB6HTICUdqdTG0phIfBzUpmqnq43XC6EHy0IY122ER/Fb3rxlG3sSYcuT4NkmLvTm1Q
4NtrlffdPAifpNWf+sQycfy0Q9FTD6yHe1PTsX0Epo4h5GlAzDZPTuTir+0YMDhcfsQEld+YHERi
vCZrQ4KyvUcp6buoUiNex/ZpcnEOibl7UExfZt62VLMDgqJ28qnYV0w4yGcpDMHV1IxtoafAvLhe
hKq54cEPA3mMZFCiPBTPnWKbu377n40qvZAuaXH5nv3ejhIxWuYgXcEXv0jPKRPxSv8mOBE8mAm4
RYpSC9Rz9HDpPGACnn5/C6yAHE3GoTmcM+ihq7NXZ5S6fj/f6Lrvj21EQzVfQfFq9n8J+OhYczEi
cc8kdDDbGAv+MWqDHvSOsBiOY5HESmLq1xSXgungMp5vzda178PYv9xj+N/i+Kz+QIbVRAd2H0hf
uTtOXugdg8/Ap6PVolFed9+6EIwLhPEVT7OjiBTVMy6qPvQTu/tuTg5s7roiS4u9dElZn35KKW2B
CVJMdiFfiDRlLZYweVtCzt0/BCb6Sf0PGml0XHRrbSMeKQ/D6/Y/uSO0bOe5kM6ZWt8yQLjiT+0x
IZLfe4VxAVHWAY5DCSfP0dg17ZsqNj9i2qVWvFFP8srpesRXDM1cRfquRFV88SphFxDOfGIm0Q2h
A5M2xeAfgLk6X/AxdsnO5FlopQUzbikD04a418PtYASKpekcpZ8N01VkFYvZvDivr8A4n2sQR2S6
lg2uYdkmyNjhmFu4b1kvcxpwaVhj/JoblbBElD3CTVK8a6K0lZxkG9hXrSo9EXIibT55+w9vXXDm
zys6fas4suaWLGxGH4RxnRcoWvDdmIOGcIQlYvC/VliU847bLlvy9xZN24x1/2Er2j1Y23772bn0
qtqBCcuBoBRoxm5XuLFtKGfct+rFRXl5BcDASHMHliuCVwvzIOHGzm2hpAs1LA+0J1JKDwr49+Lu
D17+ZcLyA1+iz6Rmx8Qvcrtwl/uLr0pYDNZx1OwL0VJagzd/Xu0R5nOe6fK1ENq4T5Kh45DKaFKB
ih0ZEfIqc+cx4eLQ9dFO9pO4EFEHiL2NeXdUrtKOPGGxlG9D944EWItbRSQWFSzmMFzLN+ETyBYY
P6Y2p6DwtYLEI3At4C8KHpKmZFEHX8Y94SlMaggNOzeLwBo73xkFD+LZu8c2YzgQs8Fyytnk5+/n
m7vsSyjdKgKZtaCGTOzlwn6RhjUKFWZDVMKIwPyn0w55bwnp3nUAQULza5k8reR/s2Iithm0VtK3
eUXK+aHvdXxk0Xp3fWXn5l6K+FTNA+eNP3uQl6wYsxS49KWbQ29xyBACZ9Tclf2N4a39l1eQjAJg
v5GtVt3v2CEnoZVvTrJer116+QfrGThpGoguh5mrHlwYdoEZNICkeky9SJydm/1n/EvEllLOyvEQ
pZ1N1LiojCKEeUiIPT/um6u2ktytpVlbTGge6GH/2oxFNCEFnfwJdRWA5mzJUK6/IEMxN/QpLEP2
xZF5uu2ZggIzVJvV+52NfydadIUR9RWEOU5fFmImxQFg83X/i4Wx+UDP/mBTH9FFKwMDATPd23zu
6a+0fCUJCcZBO32cLlonZ/3ELSDIldUnaZImkmfVjyXKv+fw5Vy3/j4023uau3bmBoJpd1+fznRP
o7xvqaH7ndn2/l1qOG7346eYRF8V1hna3OpzHMJrkMknSE8TG0aeBdwqmxqWRFheGcxIpB/Ebkv0
RO5Bgr8LS5iCeRBlzaa8apInOjYh18FYM/UybBfQkjHKFD2W0TwW+29xdwqAWolLhF2ttoxOIlnn
Z0T0HHylGoKz4XJJCu+IYolMuX8TFaeDfPu0RtnjsQNGT1Wbuntt5zLYLsTE0zlz+CJTrRJHuT7t
Mgz8zMNtGQAwgOwkWXPqwXEAUNkAVlWyziyb0i7vLilA6FJuxaI4f6TtxbzLEt39UDv5m7kpdfxV
t1twabqzB+8cayEHQER03j8zKqu0+8XHydn5k4j++jeMJdkHx/gCBMqmuFEbcseFUzKYJgwNs6h6
lIQJemvEMiVi5+M6oRfBZPVljq/eWoj7RrBCU4xKbwc07bcKSak4piLj9XG9W5gSUFMwI1ZObW7l
ur1wEeB5RSQOjb9FVX58n06gx4uPlaQ8oCiBGN3IauJxDUFJ8fWr6O9rKgZdsqiqZSWsxVut5UWL
hZVd27759IuITkFq9IU6KvDilFpEfwu7BbEMFqK40Cd2c7LPSoogoOti3JY9T+4EdgBAkAHzIrPc
iBiMeHLXC6tEwSzhNVnzqcvM2gmrTlFabUS148j+e8ES8bRq+8APPyaqMPYA1WV/V1Mx95qDbZ47
UsDWeT9RgDrX1kbj+l2hsjW7DFsheqc0K4Soof4B8p7Kh5JysFzEJhfHq2U/AWV37JdW2cY92S/X
Nk+z1Ftg90sw1vNBstCYqhm3czakqt1eUTHDAe+azx7n8KoSAbQrhZO9w0LuuIbU2lR5VgDjFWJj
MApHk7EmLiXi9IJDk5rzueYx3xkHK4M6CxHF7aTGJDWVo1c/rvWotl+HzF1BkeVBFmEhvLDMgPNl
v/GnT3zNNmsZPX+wGr2jNTXet0fM1P07hEQ9GFbdRjHSWOFVIHybaQHYxbl71RLMGOWuzuUNuCs3
utwhhU/xf/i/D+YqDNOK7yxldFw33IIG5vP1VADzrGGmA+mi+As2h/57J0frhMopJcqOivEC5kXP
FU7LtZN/IxiE7nnBKnti7gOG33F3v2d6DTlQVug7IOuybTA0/jUTOhJDX8QFrO3LgO6+sfjiIVqX
j1w0BYcIawzRW6PLRNam4VfJoAEWBgiY9gFmQHq0hW90HIu/f2uqFkWx0htTMmdfjN7C04HEE88k
wXM6OQOC5magpHsGnFsffZ/leWIU6hFEE3rb4q2ufTyNIFUqcDnOB3K+byoDEig6LTWwdFIhZ2a0
hofgA9lq3Lkttn2e2SZD/wILBRxE6Y+tea1tmw2tsqft2V/ziHVEmGmF35KNnGBfpqmvmAY3bR+y
/6L2L4d6kejLiwCc29KCTou0ScSoZmvQ7S9QmrpV6IQ+mtkfi8A/hJlM8oRgHWOf1Tt6IqcG01ks
/CU8YOeDXPU1I1+WaKqWXNFJe2MHwutjtRy2qJ29rAG2P3JevNJWB7AJ+76VCJTt09BGS15vVBOj
94rRUGo+LQkv73kl5XzgXtyAsY+yKVcUuPQQ3oWWRCZ2A5qAR6NnK5qEWn4uBYjjAspHZjoNObEK
e2DpX/s35/MI42SfwaO8QrMTu6SsMlJsxB98ZkRSsHw6Sc7Uuvv++Ra84tnbSGNwJ9fuz0G1ZPEq
2evNoOFlJdwVEAe/6P3JkMGGgwR7mvpSJ3Hm8gLuASzgyM0IZ22hf9UCyuBxTgBLbLsbxsctOI+d
yLDAQJ01sGbdWzbS+eDOdeBseawMjn21u6j+Pn5HJPSx3Hu1PaiQ1+52gT6Z7oOZ/+oQVKtC71kT
xW/0irMGOH7ckrTsUjeYdmXmCH2Ew3thu8zKXRyIaiAC08wG7+VMC6mVnxJMlNxcsvp/sHTGLfqD
l5fDLayK1SKb9pieZevmfL7QCTJIW7qO2uuyCnQFHBMkafb+5Sgr4iFD7GuQ/CGL+mlPKnCI53pc
Fgty4yOw5JJ9gomM9qxL0VoWpVxH1fN/sIRdUX+APO4zk01bmQAQDXctyStro7kU2tPq1FmzF3zh
ms0hRu8pakInSOrcs+6Xtz9V59QdT5m6OJOgjEOMH4xR9pMJEHMDe2yAgRBRxLW2lbrL1y5Tt16Z
ECfthHg+QKc8j+2tcGbwwPOOEar4XjEXoGiPrcdMcVGJylD1SvL+Q9onA2BQzICoXYRg4SMaAXBe
pwvTT/0vMjzVKrDT89dQicnqaKitir5DtTF6f4ltDZlA2stoUQ33QluE0pEsaQ44KOAhp2ZxKvIz
DXwZfLI1LkMLqxuXBHmiA0lIPB0w/ZLd9hwtEN19oa4m8kx6j2iXub3QM1XyvtikpVzmQ1ZpHE91
uXT7AL+s/30MUKCrWxR3WtdFRe2QEWRb5jR+FM/WYfKRzuLTsIkQl8elPGQN6tQpYLpRs5IU1yyC
UUgDR6mZgPEE9dbRbFCmZIJbtO7bDvv0BcbZCgdZJ3y0dQAdOtWPR3W+HGDt1wkzbEaxc6r8CgQU
M91ySMwJu8cwbxIprWXx8eaM5UkSN6rJVMmTacMjmlr7jVYHl1UMSB8rWhXXgQZlx4KPgtNIjVxF
qmOHLwoKLBoSSYRdGgExTuLxFAl2QpGqEDnWNC5s6hrzFpc1LVsAMd4bSYWepZb0u+6N6dxde4Tk
1V9cHCJQPMhgpsDrlSXmKTYM4m2zSOUjZb1Jfmgk949B1NsgyM5VSnMh7N0JVKVE+zpSocNe/NVW
vsQKXsqKZCtFvn99t7SXRIVCs43iFWcRYzRkn2uCw8rX13yfyyKjV8BzetChzMk3qZlpF7kGuReU
84DmyLFbb4qTYSZyAkujkDrl8GtKi+5Ig+ujQq3lchwUY7xyLEcJD+S2Ah0pihYDUClBercxToJT
S6wuUd0C5T8DAuMKYKns3Ul/rie61w4arjQ9KJO4+Uv0ejPGTyjg4vJJ6jFUVvVOsX8mFRSCDPbC
E06WMXS+kV2SRGyYmNpsOiG+0CppJbX2UBg7wAljdXTkruOWAznkS+cP1NWdvvmmTJQ19yFsC1ts
1sbdfhnD0+p/S8FCemR0LPvwmdoIcMVuxXurq4Ht/LvS238kcpxn3kqgHAZqRoHie7TlhFgr5crt
rQNd8hebjY0fHdFfA/jvj2c8ZDgaKp4Quymvnc+Hso6CD6wyY7K3CE/N7Ba4B4e0JTRewm6+imEN
v63qBXphlgapVzO80nTaz2jG2fDJoyU1+njypkWbATbrwrucNWAkTdkG6nlZpoHoyuKhmPrbxrPr
DqRiwEefQC329vDcZu6I8XrZk0R3hrNnVhia72ap5QFPEI9Td0e9DS2mklHC9OhAt4BpHFXipvYU
I4KOw0v8n98Pf5s5psbAPOQwKI6KbJEG7kdoJcgGOzlhZZavsJN68nX/khmDBWXybJni5MHWoibQ
55CPvQbjJs4lNc0HeI8Lm1UsPr17prOfNnsT3bfiLv3dNVAjkixiGs2VAvuNq2nfohy5EIDOfgfh
vBmlt8LkFiWf5s2xWmkdeVp4BL72ojfhVVfPkkWCaO9KeyKA0pURo12TDtxJ4iCw8znrgeJsVdRq
FIfmRipdnmdj1ybzeANx2YARyex+IZCLUD5W56WjzDwLg+eBhzaggodSa8WKgqZzNe0mtPjuBif9
aE4eztIcbeVUFr+fa3VHHgTEQs4hhV9SvKj9jT7TmBjM7oYyF6+RENnLlB4oAIADrPzU3PwJDQ7Q
KHCfp+4BjFsBOFXWZ6Ho7ShoK+INn+hO062FZS7atq7BtiYxqfHeB7htBfR0J9D6OEi/QhzhdwLl
Zh8x829hRp7n6wC+7QFMpEJMvRuhkeBEtX1ssKt9J4MF5+wbCAGnygx0h5FoHPQhx1RaIS5Cu3P/
tK/B0BfC66A5ziE3lKd/SoYkBic1bLaWzcFAIYaqbfp+RP8aZ4n2k3LtCZ/6tta8KbUziLmBJ1fm
HjS1ZHSxa0CQwwVrGSVxRZ3XVt+CqoLVlUScXH+mfEd0WCZ5HNE3cMzQOY5QCJBJYgFLs8sVMsHD
sKBkTQVzpmqjFZ+ns6k9LbQAkax0Py7tpOuZ++dXi9nfxMy6+i1b6qKSFsIV6tEnka/Xofdd4mMP
LjwBVFq3Y56bgD+WmCxvpNArXbs3vn7KPJq8PLR8PVun61HIUpYtbGT9D8SN0x1uupJyvHrFfqCa
x/Td7uSowxSFHxVe29GtWsPyZ4UNDZ9svg1m/4V+InqJ/NwVyqFSlSAZZ9Oc9oCFeo24C0tHigqx
LTQdREoceagmh0pMficrXwYMmJxlF51m9iGMvs5p1j6smL2sD1w8cT+Ng5Xtyz9I5fFNWgtLKwGd
669R0vMfgkUyLS/ubvtgluBHgupNFj60zlILMDxZh51MmpoFJkHZIzoyZLtYmQxRKbwMIAPLmqRn
zSgp7vy7KKvSwtSMYP+dWo/I0jjXVsQ0Z7XdtAsiPZ8StqJesoKUF1tYdgzaJ9f9FR5dd0F5cTdx
nN09rSLv5UOIPOWMZrsxpygRnxenPjLV2FDSGySpzoh9mrfIkhzBAtb+JTY99OhOhOYbVKBgNlL0
0vrT+QC5MQBZewIm3GGk+OntCoz/QTqiH7tkmJdTufI3Ygw3B8wlcJRYR+kX1JFAnYT2EYp4J2xx
qL5jMkFObjgcDj3kprZESVTeT/IHDgTg1lHnYjjsvobCEhyXl99IVwiMMhKGdcJWRNQFAj+8jrLc
PUj9unmqc8fSta7ZGR5cDqlTm+skB0uqz6GEUoKH+E/X+A2wXp/9Pk7p4ISI8gqr4bXu1iJ7V2l4
e/Ah7t7Jw3pnBDvxaiKiVSjI/8ewYWvhZ5sbrDd/3yKqMwDe2TG2DQ48yPT2Dw081pyHcEzT1FNJ
OeeOp+x5KWCTvG5jUY+FPEE2c57FeHw8RYMwiPg7Rxq7urb26mPf75SN37OGHOP8fzG1bz6VhbMJ
oahdIKj3dKcj28gmYlTEJBTq0xVnMVZzgBE3aOPzT5yqx4+DzuPkSmzYUQeo74fCHmUjf7aYv8A2
MmpwUTsud/VCPQRhzX7NEgd3OWm7kvLUwyM5lTcvNVsvMM8gK4Fj5uTMR1ht5KTF4dGcjVUmduQH
4fxQiKofZPFRoCq89vQD3QexxIHcnqKKT5l4FGJME2TukT+TJe2mKN817JS0+6xBdkMnNNok2nEe
llO5FaBAAQI4UcSjr+WrnAoofMI5f5mgt6HmMFe7HAfhDs3knMKEGzq60qtZiEi3oQ9a8LhMDD6x
lgLFp7Au6VkgkxoYW25ICA206BvZPYnyV5f91Z2cXqMXNxWk5VQzrnrpPR+0HSdY7PaPD6u9yBbz
7XWbIxYkmRdwyD1b/TyatX8MrWSd8r0DgetmgcTydxqPqPObEqgLO4s3TSAqjfd6raI9FnhszkR/
f2CM+/JgqQIBDxV0iTHCJ49vegyFiyHQuHJj66eO/4a/UkLRWxFclUNNS2/Q3F9yiY5ikA7t1mGT
m/y+TwX/ovkcwRD+Y/vHPdRK/UmM0tDgJdqQUIkIpnRLNmvm6ZOk9tFIZxroFb7lZa2+YpiXGUGv
C84y0ioDxnkZ+uccb506XrhXska8dDzK0nXNqHxNzY6EzEet7fC20YvqHcrKkgnSsmQ3otnrtxmt
W17CXPGZxBDbKcq/5xLRjSgiTmjDf9zPH+fgKlrnesMO7hWhf6xHmfCZw7CEmuGvHa8/ni1CtfYk
CVIWlE1VP6gKVdeia6Zboczbo1DkoY3YhjyGeDoUIzrX73wqfoO4GG2H+8cSDH8uyL7nm9rQe39V
6ge46BuLGz4AmAdPR3YFsrFdBvARBCauD0iwHQiliq18kY5KfacYioHNgI7WFPPbMd32bR6i+gBo
agk9BrvDjZFfOdK/nKp+pNk6AtZtwcx8Z0d0VBjW1v2XVSJ1NnUMMB2QaTzbrP6e5++UmdNR/h7T
mCKJZs23hjP8WLHAr+oa+5oBKdum7ePdFsfWGkeRDtZE+LB+QIiOj2N6cCWgV1VLw4/TSnwQYBcL
svfsOpxZzM/5IjIqWrrewa76cvhWm6Kx//Rxo7fnGICp0tvvvcL2Xn/lMMzailEHYCIObSeY0UKK
Z/V3o6Ow+CaWU+qmC9SMh6f5qZZxlvG8j0gocHrhIbjtfluzX8dqoUtPfXfEcilxlC4Vb1kjFrvw
m/UJKhVnmkFjSe/IFpO5HPR7Zfj66E5LQCAiS4IF01zwhixanVC5P61HnO9ImcjRC1ReaXtOzgId
orfa6TF36ZeUSD0BHBhRwFR4engO7MrmdR/tsIC9pAJfCU6u+lP2HbO5+gv2lpqSUyH9oD3HRTYd
Nl1Ra7oZZS92pkf21J5faOQK7lm+mcxif3CZ6Xp5JWxhdN+OisJ1DUm2GWPr8nDs3d2Ofw+cDhzY
yoYF4SZjwel8t6gEd9bauxePRXsS8uRVBAeuLZEQSS9pyQaALoRU44asd+/YG6lTquT9/3EDj5Jr
SX9cPM7BYn7ltO5Cv+s9k7M0r/sQULBXVxi8TSOqbmEO3HqGoiRkKaz4Q0kAs0M5e9YchOOJ6EKm
ns+BjujxQVbRJHF52zyz/tV0LNawmLMv6nVbW6gaTfderxUfRzMQad14meXyK3hyTAVklZCbd/uk
cNy+TZtFWxwUYDZP7dD58V2zIjd6jufXSZTdMGn6tUXnPf3aNmaCu+ZU9VC/HvJIJw/6JM5mt8ma
IQTX/xN+JDrUI3KIQ6bqEnhdfQIFtKBdY6FhUqSzhKqmnsPgv9qou7oumC7T2VJdZXTJoea258JN
nYln485/eloFknYATH31p12H8chOMVkRccMtBeskDo6tWgcQEaSVtJtYLvvZF8c4AeCjgR7bg8EG
F2v1OhKcR9FCS9WqRQPambbCmRQpmvgNd6bjqCt6f/OHTsAQWktmDmmLIWbU4aI6deXpSDCUovNM
t1R68BHbfs5WcGLQ+xomD3zWtd9hswCUpBGxYq+dTiY1Eq0L/Cv/SJWlCzve5zxFcb8gXz1DXM+u
pgm2f1sX5eXNS0LPBi4r+XI17rRku9qa+/suN0tQ3YtwtYCY83VjmefBu795cLeq2IKn1gCJLELR
rxi9jQCUlC5KBbcQtmysVh97giyympQezOG/tGycqbLhfETNN7C8QBhphQOkBqQnrqC76uONnmde
dK0Zp5i4GVhx90QSKgHYqNRW1917YvF3ZogZGdKAXRSKrQ+6H7qVZN6rV7piGNd5ukYI5TYzi1Pa
M2SytpKkZ3Dc6s5GFtPUTbr4YekS/ZsTo2RiaJLdu1MXXN8V1u8fCl3/feZYyrVjLCqrvoXH36wo
KSpWUd7CetFOM5b7Q3TDNvveXE76fL8mTbl8AdOpt+soPUedCtri1XmfXDwrsodNlJEFXkivemvz
qtQ2v0JpsGbiP/Vy2KCVJuhQfd1/jkLbfT9Z7wWnLNWKelAhlMhZnH76nH6Mom2XylJ2QnUBYGrw
xj2toOEE3HxJw0sTCseN4pFthJyyF/bf6h5kLdFstlcqJzBaaz0U4TLPRrjTPer1QMT/hHkXUNUh
utaXZ5n3N+OWNJEVlmxD1hrHOZ+2ue81MWgOaf8CcV7EUxpRbwqqk95VjXR0MuvNBx2hjVVuMEXp
UXF5gvBc8X6WlLv95AfAsxveuBSj7/Al5nLr71kywn1ccEhYgJ5VKEldrsv9ZE6IbknyHfIM69CC
17f6kUcSNIq2yEk5l5fbZyoPKYQYcECbbJXsGCW5mWEP9K2LxFCI2xlILFVfoXAT58xMMVqb5shY
WFVntDlUUO3Yk7Co41EF3LrqmaRPxHLpWdlnqkirM1WuKjo5zdZcKPdAV9cIxfFnrtJu+TIV7bEd
1QFqn0b5corcUGar6JxseS8rNkC9OgZazVHwe3TyQu4lXGnuRlBSksWZX8oUUz8x0XG+n8kxZuHH
NTBBmgcROVVmRocxCE2gaUFfyE6gbUvCCK/W8wquJEcKXHA648Wta8kYJxtGs8C4kcgUyQei/DII
ad6m+pxfVhIduChptgGrd5/V3ddzhLM15uSatqy8buz+Grr1LEqGMVDtEcLcDCE6NX6+gAZTNcBY
1jX63cBcPrIrrGFS/vbLkk3EbKSkq68PaHggU/rQ0Kwri5avvjPG/watTUl/aUu2uEIAIhyOq0aU
x5XAZ+Fwhj3vJbWnHlsjpePbyqwHjoiZSlX9zcpUXEqMgapDTm9t7+Ft73pH6Wh92dzEmNA5hlDD
Jp1ldRf3BhXBgYiKD9ExnbgAQcX5853s+u93o3VAOXoORumHjrogfR/UTqEk1EYMnOmuuxQVLajX
Nubx8lHiV6Wt4nQyv7RMbu/Iklw7K/kuJ449FvgGrSoazyRYIcG9UrTjm448xI/7kZO37iA4ky3z
Q48bvnvIYPTbyrO5AMpquapk1+Cd8+XLAcGP/k0TeFqIANbDJMPofcbRCHhddCFszSaM+TllKwYc
t+x2hLd3GXglpnGxfngUIizORk+grw/+jJkAJ3hhzjWNmV58jMamY7NgPBDTjhzmfMoYULMII1kI
1kBfyUh5kMI0EReu00eTOGmnyXwyAvdjGQGZcP10o2RTcNsrxIw0F8/oJyqQ6hTiNiGgLN77FBo+
gnpBUHiHHQyeOkhJ+Xm7FXlBsqgAu5zHI3JXXlSTr1+AlyQ3wJWnQ3kXRUCGg9Zgm8mj9JBpVdzI
DjK9cyxjLuYQ9rQ0t5dU9lYbpfokmBeJl4Re1A2Iqihvx7UjYiLLrhcKWWqNQP8Yv7wV5+NwAfPh
Qd4k5LsAWuk34YturnhNZlNRutjrZ9cqx/W8IYN21n4wiFXx2/TmB7Z/6AS4vhUe5OUjnhPMPhcR
LqCAEURC+ctEz4Mw0SD+hgGwHVyvhfsDg8VP+zYZi8jiHPcSvUtnGzDBa7O1pJFUKOU27/nzp8ZO
P/mo+n3Im1RvA9YRMk+78e95X/Rj54JgYESCIi7JueeG3lJ+MRMF54jSKDWzdE80WOdSj4339tgt
VgBJiJdlC0HwBDW+xndvIbOhSOACXFFWI6jX8kjzGYbxntyqKzLCmEw6pOPt8H6sOr4m3ruwRV5h
iWl3H4k2iBxUQMT5zfO1zh6MGK/bYdxYch5bQ1Pti9SmIl7p5zgf3+4/B8x8H0GWroHB5vCN+AsD
zazg1TsFCuDTjeH0s6TTKyKz5ODZALrR04vqPKN8yWLXxXR0zbhgsAeMqkzlABTgDd7ZvrFlSNKn
slQAQPFonqqtM0YMkSp52DTbRJmsLkuKHB+hyNxFCVxG/goUlkSK9hSKYSp5YQvEhDVjCGB3EZIc
jzCJe8b4MURL+DruyghbU+X3XtBuuG8761hbBKG1UYRLA+hGh+OYTzvUB44YGFs1x0J/T2sOm+T7
6Gbtd7oVqzYKMkP73zaREzZRpzfO0wFRIZQgYL61Pc5NZQ4xoxMFwMGKstD5zfdbyjXtoQqeE+2j
WKKpEqlK4T8ZLBa/8ZWuKhlzZQVHnBwkHxB2qr28d1H7ju1fddVqyH7GHHr1U4fkSVaH9t1aE3Ho
KDU9c4DB0jsQas4loE6zLn6i9VSCoIQ1LVxugDebPoDHY6r2esS5rntxB4bI8kLk2x4cYgnhAdED
IH7sJVchXLR4BodXmbA7OpfBMh4aoEhYH2/C4SZqhgjqlM+xJlYjp7GCPBcz/xjloSnaHauHghp4
Nfw0DBzwttgvRcHCqp+3kX5u45bp5OolFc+ZQJ6/6vpFzYtkBFAUj9v8GwcJMpLbiZo/ihrHndwv
MzTdpuglzGcb35dzXTH4CK0nfP/YgIyYcLddwWHgQR6fPb9Q0v6cxmeshKoyLUpIanp9KlAUas4+
+CKE86NPRX5GGmCYhCT5eWzhHnhAvW93YY1RA2wEx8NRa05P+Z6PxoeQ4kQqdKvrUlGAUvGmbfov
x8JFIIpwBRFqtZSUX+GeZio/DuTd5t0belaCGnOsPidBbU63SptvmfuHpc0BKelMhRMSh57UWaQh
va9aLo7D6Wp2HNPxs1SoyTmDURsg6K/Ff3dtI2hHrrLvHKVR06IH7OusAaBXp3+YLLhHZ1KaiHCv
lPJAd+Rz/aKDlVs6Bjy58w+Nsp8nT+G6OBbG/xKTJ3mJPosBZxLAXz1CuxscJcHczJloPRfH65sg
aIA1An/z1mwi7279KIue1lkGWFZk8NOu2m8q/cQwOKG9FR2IS7aN7FxKBI/JaveQVQ6D8VaKYyRC
Acjq938HAUaWlk8RiNb9Z8He3raAUIEWRxOQVPkjxLpwVsu2Ej1YXZkUEtaLHiwV16jWMLNIcMjv
TLFxmBFfegIipRzGIpNhgnAqpv5PFQsXFR5asKNaqandx20CCZe2aBjE0w7ArP9NaojK31VP6cA7
lLEmij4q7msbeQuSTOyNt/e8R2Ma03nXqhmhj1N1HhCTjHLt9jT6DrAsGD5DATvmgT0qjAHG9xJ/
PXczvSeDyqtaiXrzHG0t85eVLY0DnIBDas2VQ6l6drKtVVLaCN8RFavg6hxEVIxR2/suSrpYfftL
+nJq8RGIh67VeUj1ePfVy13/XOOa9L9EJFwhGTq+O75gXSBi6RAkuTV5sCHh7XAAUbL1XfNgCy6R
Ta5gBAed6VC+9fpY30BhiILmi5A9PUVOmjCU9gUptiqprYjND/R5e0bNIbR5zBc4M+ZPRY26nKYU
ippfqvOI4ZlI6jw/0K3uUGawJCqduvSByy1MfrC5vtOLqEBwM3Vilxg+vEfsfmnVSh7nZQ1O5j4D
/xWhHEAt+FgDhbqFVzgaA4vyFvMNjP4GV4oLQtTv3rIVPPoJFMpLp1dGdIs6i8Yu/X8bCF2dYFjy
Pt1S5O4jwCJtLA8AnfOjzTcl6qysjtM/bQCBK1T/QwJEUBX4E1YLNp6sBAiIYs4DZ2pzxcpsSok0
fytLhN+MH5qjW4XAwMmUJP4cjLgnUW8ONxDVQdz1RMNKpQb1ctPmfEHTKn/mExeEHZqxnFdkkpoJ
BjdQ8bb4nIm3gBgRXN4dpaiQAGFtT/wgNQ1vP0ES0uAIVMRMHsdkU2KhdPP94KdqAO47gYPU5E1p
7Q54UrXoIyrdWWYlIRLzIDtBjBY+DhECzcS1+8HeMUN89GVBf2c0renYSw3tNn+Xb6kK7pqRydzZ
qaA+4m/z3KcTFnz++WQw77p6z1IUKTg4J8attVbeTdKbtgOer5TORAeD6AI6Ab3GEn8aqHvYjq5f
bROvJ0o8KDS/YguPzNLDqpIKjybGwIO++yH/VfRYPxk/Az5bKaUbPN/lUoADgeJd7y6G89Kl5y/L
inxVGXT9BS/pv/dWYbXxNc39aybwIzKx6I2bH2U3NJ8Ugs4nUTqn7hEmQV5TZ6242WdHlrVbMGYJ
dmI/sc50cCmtSJq3W5vUP8Q9AADwPGIeL0NTnGLiNNzdYNLci9V1dR0bRnynQvDNH6Zmvm3NzeTi
khF6YStDQ/I7L1teYpwllydJdS4nf6VRyI9efNf9K44aqjSobOUxeFRMNK33yWazYjoDitgFg1I2
Js61rrgCuMmAQ0VtUpOQcZI95PSfKEsYJh8W6kmOMEqiatIXQpdW1J9vdhx+q2sbL7nTp1+lds0F
aNk6HDB9EkVvuvoDXhM46QtFaM2RcsfwI7XYcwkJdIIYiK+UIf7oWgYl79tyvhaAel3RaLQ2v6cx
Kk7mTD52hO3+uiTL5mNDG/e6VEFR3G5/rhlEjieqn2cAprtsxrjgqt6/BCSnCyVsAyjvKVWCdzTg
v70Sk+irGV4UXUT5V3pxiKN1mF6eJpyyRhTIFUU2CjsAl1T5LKCvEykbMRAz/sE++N/JhqliC7j2
Bdf4wC94CjBFYA2bgjIFo7i8fdG2/mqaRQglgnro2KBgYw5yA3j9ce1rUvUtp+bC/U/kbSgwzu+o
2x1Sc1V5R4NmWhL9WXWf7e8jW9+6bVxxQodQ2UcmFli6/NPHuieFS7fPTKzOTzuBhncscQqnMDZs
5A7YXZk4uw5PZK7WK+CThort8hIT9TtNiVyiFBpjmjBtuI7gFf61NB0PiQvuUg0rOmkc4GAdTvgP
sI9V9pbpIXTNXNZKbBuxpme+wEbAMxMorqBVZT3i4SIdoPDLC+aK0MX74hJyBN8ejZEt6GqQcHas
ws5SPouPRfNx7805bjJfpeCyTrBtiwLEytPi8AS0A3gjIDoat453iPbme1vQKh8fQyxwNVXTdnyo
nCbdhTIU/yF/9lJjXGWTglJkOhdd5cuCIply06RihPS5hY8vbzISMgaA9bW/xTD+vszskxcCkz1+
j1DuIb08G/gxWUNKYx1uX00Y4Ih50R+52Gg6arpnYbfb/9VPFQCG49h0ZI8cBmif2jOEtZuXy2lu
aNPtkjEe5X2vCgf4eMlMU39oDdYqsUUmE1dy1D6dl65T8TeBnLIOUsh7dUKBHBGyXzX0xHQGJVe1
iii0qsnK8RdTEbGfvO38r/NuxU85SPZqqSZl4FhCe+uj5DB4xC1COBTi+juw3X1TibIAbMUNUAIa
2sbRv4rAMc33JhyJSZnga6B4TGDCMbfZbqEg2SFzhZM1IevhepM22TW7IU55VV6hAebXAdmC3YKo
kKTUaS7e7jBBQ49eAHzLToXS0yVTEC88Uic385XvS9FbooeZfN9sohge43E8kIJaHCqii25qdviY
ii7FGwvsR+olEXI2m58dwNUnF3SfdPfAYl+mraoqb6u9zDaJbKk73D9TOAybR1JREvxeSpbajT9f
Q3UGeLOTXeU/gCmpxAyHbaBnIrp4/+lwt1NRAH+sXSbV0E5eEGyjYuXhN7oms7//e5xQnd4oqpe7
i1S9fMj19YLpER4WvCySY+/r3vtuaz41MgbLpdCYXcg2mDycehlwHR4VNrpGCV8oh6uGwszpHB+t
l3WLYxOcsJtzXzMHk8T6Oiaa0r2mVP7Bymi4OtJ3zz+Agdby72Rk1A78Cn0WPpLwCyit63LW43ti
BD8DYScyuFYh8CeiX+QBWGAqBJbsW+EohpNgRxYm1OvLAHWWa68kTfKgayFR5i0j6IRbSRv7m9NA
vJBQVo/EhRoKQLWKyJXgyYCDt3zdGHzIfzirF3xNvdQqh3Fwnzv7ywS1Ug7h8fThF6Fq+OFVYIPw
l8BviEPiz2FZ+obU9MEGnVYhGTEyJbI1nO3X8LruR5TXtGf6FFBS7FUwdr+/5RWrXhaIBxgJ7cnb
GlrqGxrvrXykkxP9zan8WLGbpGPN2BnnudxVLltSMPykxr7YDZNuv6S1IWnJlzHbFhFsehu1scUx
G7ViN4TeuGbODnREusTEaQzQZ9rTJu2KAO6t7kDZOJyD4IA+gEoq7c0i7txIFPQkZlng6/itDLcM
t3pNpgvtOb0tesHTGGyrDPxQuMnbH39JHIPYUWfB6j7mkPV/CKmHifcaln8Mvi1RiKdlnt7Eydu8
3Hs3pcCrsASM5a8TObNlVkkdBi7j7gKEFmqKsmmqs/PsuRC+gNqwtuG3TxTddp4qFnOFdQkrp8kV
6XqZLYCbRnD2Pnr9R/YsGUgwHRr9qWN2bfkDEMbAUmVYnSz8B8onKXfGeexK0a3sVLZ9O20Ete2z
7M5fatBEL+M1e0uJfBQokhFFmmDtd11EEKjzWOQAgeKSlGM04RAo5fbLHUpBFDwiw47h0kD81Jea
X7G6vVY9Tq6aYfZJ8YOXo0ZQ26WuM8Vq7frxC+X+EF+aqtE9EhRGEzIocs4gsV3uj0A6ydH6u3xS
asj0zp9pTRJDjMvPuj6D6uAWW1oH0RMLTfboG6wktbJcia2L4gsaza2hhCkzOuPaV5ZKXtYBOgby
R1rtXjI3vmlBd38Zyqfz4X+zoZo1K9WJ4dxKEvzjyi59YbxMpIJivRewzm4/jSz+d/ls+dkf5CLM
Xe6WE707zfeRuvn1byJgXefvkbmYygnmKa4so31c2nKmuWzf/qGPpbuEboYPTmckALW3YPQKL+xZ
vvxMzjBYfa9cs/6yWwUBbUPiW/s1rg0pXoFvOJXq90ksXfw523pnJUJPdBqdmEgmEBu9vlXzpYef
PBKt8M/9U+LYbrdZQ8Ox0NfV69wkVsh5IL4GTiPIdcj8e0lleNFhcNOvQVIfm4NFn22cXIrAdoYm
lttlDjetdPxO/Tnzl1AvPb0HYGJU0yl9G/zYc7F/JGJWB+J9k2OoW7AykEjeUgjo9lf1eT8glRnW
d8qkjzHs2fJrqdEn+0MRsvwyos+IIP6wJNdLfsOhn69dPFNwDHid2IV3eyaOoIZGu+jDoUfusSX+
wFoXQ+wSF/RHzSZtJ4aIJmU5U44ahIa2AIEjVb6rZJ32Hiic8QE07ts+PY35q4Uot9kzJOj28IhK
InnX0XcyRJ3viG/p8vyRSHH6/G2+wGYI9TSV//n9CMKD+QlA/QyvA/HrO0aicmW1B2t2QeRWuL6S
S2qxHiNX58Hkp485pLqe711WgTbLfaLFsPWQ1PIjUdnjLrjWhWudZoSPifc/KgWip5VdZ4S+Jml6
PApfWMYv4UuQcMe7oHalO55qlLTyX7ES5DSyAbXthBRQHV72yTv0/caesGV98STyJLVKdRk3w3r3
lmsyXuX3ltMgz4wSkshksKdDfAUtjEAodiUm2q6kjXaYfWkZBfc7AfjlIj5FV87M22fN6jYoj6RL
ai3o0C/He9xhQjIrh8XnaIJswGP4BoOnUELnDjt7oIsSevOUCeESj+eIByU8th1aCeXlot76HyMr
0i+dynit/hl6cfEd07iCkqu3//GtFps8DtgZMwM+DGmwAB3g0eL1AJbU4ljoOnl8yD8r7QrRVkRN
HV14jyq0ZstkMpLu/HcbSL2Ph8t0qbgN1rgMPLR+FRCyubSzxPz3tiLHZC3xcxkZZ9BNa/SWuKAx
aj0HmYkIztcSpHjMe6zUHrRUza+tdJFR7LmmXuhHrTBIPyn0En2Fm6AT5okaiRlRRQZNu95o+biu
bEkMlFSecBekL5vV+omfxPeX8+9tzghHptZHTOL5qVLGkDCpb39B6aBLJSFSfJ1QEM1gzc0XZ8oj
gkj4zB4zp7YDRq7YpQ9rAduGyueZe2mUibAdgKW0Cscos6XFcnU4dl8hgwM+33QlcOMoLMe4+aUy
3P+wL8kkidbUz0FwRtfwrlcOkv8NpF97pvFN6cM/Q9yue8TvwOguGA94v0JdHntOdjaAsEL6238M
BmtrM7jlrUC4fS8w4IhMYfnMu/EiwwdjPqBc4nxi04EjEm7te49NPOG863g1MDu+iQgOt9yUa9UR
wK982aBiyH5SSpTr6xYzB2FlNRmeEMNyLcUmrLh/sdVQ5GipmByr/Ha1Ia4Naw8XQ8zSX1k7a77I
QWPWUd9OX5KAkcmipUfsUssHkHhzOs4uio5Tts3Hfz1S4GkAK39XsBTb4uOtMwpKo7NMoFYgbTLB
CQwkcyhKQS7Y5s1STUkKATs/Q2RhK7+vMDufMIH6eW70OgIglsP0wfJ7UVCMbYOhKQZktHAaelP9
8hUaGJJds3gFj+G3lcX0iy8EhR6Jn0BmpymJKDJyCvEEfcf7r7qoywDNsPtzPVYMvFRjQkLkGiAT
HjcspKFOExmhAWLLeLyR6qVFIvBKjXQ9bOA/RJq5ChzsdeONJvPfVwKvDz2u+fRNvvo6SXaCdSwH
UX6V5sFSEqs/b5RqK63RykrYs9HBIoikPkhaFYbgXk72pYt715WUcDpBuqmOQhs/WY9QTWfkAMwj
bAhUF9CfnUDa0W1ihOmLoSoDWRvEM455a+9xAmqlRiyCREH7UvsK2EsAu5Ti9narRso0v58aWQJ5
cYshPiTS1hZNDtj5r+S3Fhy4DwtPJ0+dzNSb7YyPFz0Y4CUX0+VqN3Iy73w1354X2j/syB8JzPXy
nB8ikyVAD2Y2c0x318gV/A6FJQGd85H40LYZfewFLHvTIxn+H7zYzSkPEroAS6PIsPQk2hlwcz15
36YBM/meW6Qpcl+qxtd9cNTtbcnRZ1gM4I7vV3fz1cpq2LW/a5r7deLDQwPBCfYzBev8E1euJr97
eptX/4KgrbGeddSuuovWrSBBpc6r4ob7ipMstZdnHvRCP8Vcmwir4CfWzjNmdV0DWn1uv7sntTWQ
EJ5XtvdhueFWcMLg8/1s3q7LWTU6Y0qIeP+h/pxE9/SIxl6XjOip9+Wsmcr6ZJF8STLD+31/hPiy
+LXFbmMQr/x3tQh0pNfuyI+4Ak00tTkwxUhhPYM49HkYmsxtg3qGBHAB666E/c4TPA19RgHi92xE
hrOyi8+9/6qSArWPRXJsfeleU+i8hOXqSN7O16CUr3AjMhF0I+2F21PmNEH6RcF3ffdW+FW6jRKk
3Jadh4iYoeff9AJx9QNqZQC3ZtaN0bd+xGzyV3R+bAILT8+veM0B0hgiH5sQzaRL21kl8EYXF87v
dPYFH5DUjThnqECwJwhwgCS/Qv1LPwKfgEvZhTeSxtQGcpBGNXQxqEIra7wBvvFX+mDBL3Z8e8IW
eFtAshAeqkXAiFioOXlzMT49k99bPegjESHKiSyrP9D11qlujy9Y4rS5Gx0DMMkn12W8m51vFCvm
JnhkxKKSeoJ9ZxgXawenfLg52zJkMI1LHayiVHh5xX7tDKAVrn2fncqzlIto9DhQOWEP8aYlBNaR
H4cK0qLuMinv73BG5GqXWJhxMcSuKz9Y/h0kS+O0+CituAddlP8PHgAsnkFJMZVAEZEVxu0evZ0F
ga60HOQpHvsx8W3diLZRgDybWwX3buIei16vrmD9o6S3dGRQvU+GabMy8U04vXoU47w9GFuRKVpn
aaxZVjE2heXWtxZ6EqdfB3XrP03GkfsARW+HZKENARGbOViT5BHryRF5npt20uc9iNT23D2MH2g5
U1K+6uFVTQKHZkBKt6pJXXIbRVtqOGXZ2yQnWwiGxkz9j1THQJ7VuGgWfuLyW5EmJvNHidbCb8Fk
IqBI4RQtwe5kLWZotp5HI4OWkt1ImWyk4BeJNYthzJyCeCji8A/3vYXDfxKvlZV36teagDLHB1wC
yhLshlda9s4bwT56krMy/mHXboBt9LcgHxmDavcCEw7bzjDxNUixou6+Q9KEZdI/THFeXmiUTYXO
3nzZobVn3/l1lI1S9vwbS3IKL7wud2945Pb8xvm4JjxMONLzNKPc2+3nPk2cujGJt8/wtMeAAZWv
eKRNM/SwAxeGM5cLVKA3sZ59xMXHDyvMFmoKy1bO61ORf9t1adoMm1bidqlciDchmi/ggriP9OkP
LxSTRczYevHvOzFWAYwxh0gxX2WnJdSDV1s8KL645yQMGX1FlnZK+93/7v1GEtwzQY1qAY5ZGhHn
1s0O3oPg3uecXNaRylkb5a2nNn5aAml79kNoQLkLeuXADLJPm2wlPsYQqjJgBusk3N+MttHkboWI
/Ij9BiOOlCXwfLucdskj6wRBOdHm13Haz8hIHTaoafbAgrVGZM33juuh4t1HxcVgr9vuUsAqF8Ho
rFod3gRkxgp7N52TgckAiWUnq7ZOToUq6gvA172dH0eS3S/7nRdtAosGxfEgkiJKocnxJpkAEqeb
BnJDOhqpd2xZNR3WlrLql6HxSeHlZLvg7coUJwIFLF2QkC0WXD9clGSA1wG8uoGzcP7oUcEx6XBL
g6J6cuERsHcSK4optWax0xZUXFhFMLp7W/UAyUy7Q46jFdL7GZURmw2yh1PNPERNc/yRUGMC+Fkb
53uNMb69AT40VNedEtBq27d7SRU4SbyO9LjSj1t76hZ3QkNCecCgrxr8IGboh8qDmOaQgqdpw5aY
AXrt6gln6DHjbxx4BpNIf95exEEHN16CQvpobarZwsZn7jkDdy3UOc2FZJsAffjGMz71nMTYF99H
dP/IqLfgl5u/fvayUQClJHaDgk690HP4kCEa6xbSpUz4HOUp+9uuitNo+95jx0MRDI6fUvfqmgKF
o5yFLFBuTa7HgvLqL+TBPBWJUmz/ipHGaXMDLPXGEI6VqieH4/ztejPqOkDbCg3ryycqMeKFG56O
M5ScKEHCwP8nXqWjdXp6u3YNhvwQp9nQtw7kvff6gOtpNJrV/FpA6LlHLiSlm/dPxuOuQqXOk6Lh
xofLHPwp5LSN+ofTv5/HUfiRpQI3z2bTKJZoAOJ4JGLD7tffqr4BPyQ55Lydufsdcc/ZVuMl3W/l
rlePjxRrhQ/4IZ95ucXFa2J81xTiv69ch5pFroBRbJucEQz8uU+Axzwp8BKo6Wc/kaewhnKM57TZ
87Rfx6mOTtuKLvhreK/Getb8wFAJf8MZwSystgHlp8BNdL9O6W8ZhVJcfEGOAhxEF3xLWPFB1+Lk
0FT4KT+t4415MQu74nJuyTIPAhHE7r90V6Alfhk7CRTrLlh5zYyiS3gpncuwKGgjJ2t+GvDXirNI
B04yIAyFf278MZhwatfZaE1iOMS8vYBHRH9Vwe0PYDOTlVzwbdoj+DCRoiQ5uXNFfmgAzLCkwMtH
pI9kjAzXcy30eHnr/W5ar5cKJ8A7f5t4VJcslVqno9aUt6+rwWMBpio+t+6aJCuM5IXFVJSVq5vu
EvY7CN9Bl4rZYgc/86EeQYM/kfbtLmmJ5zMuNVudzeeLFcg/x2c4NDuXQ9Yvp2/fv26Msp0f1LSM
sit1h5Snq5qVgnrus40HbA2CaWncvdzqI/vllnrp3t/45nOqL/JPjONyDfOWtRD2wXifqJKAONfn
cpgr+udgx5NsXUuDzESoOz+z70zGVWQHRV7AG1NwXOvic0Iccs/35k53WM9oGac+Th1BE5carnfn
aXYXQvyJ6xLg+94GQ92gTKhCu/HVpemNyd2B4zcxZTQijZR0+dLDO7+gp5wGEryMPPNCiOjH8eDI
b/LyRZdgDM448DnbUdRSBB8LKJAYKDZwqTLvRX3mpavSXeFkis+sprL9Nn22HvYHUjTPTNpydNy2
ac1kptJsJ1VtJViX/971C+UyRYEWebaDo/bSmvFOAriLlzy7AFeqOPd3CVww5IeIT0Lbk1XJ1zmL
AlQb9dC0VO7/2shu77lbJwoi1SLUkfZ70+0RjXI4tJLNgh0NWzL+4jsgfPLP4WrOx/0e8NB0ta9M
whqTdvfO/uDCk65qScnl0Cb/cnOc7wLyvmVYr/lKVcGJYhAFI0i5r/ul4LcY11UNNxSy5iUGXq2G
d17L2Z3HbjkyoIDLQiOt69/hwe8TszQlaMkAH6Rkv1RTXLqeMD0ZaB4ZWhFTGfP2BSGkTlDayY91
NvP9RVq31j4XMKrmTga1YVbGX8h+mgsoNxSaDaPbSx+mBUOGxjuXw6RDQr+0SXJX3gOiMWsPizhE
mySvlEYlD6eL9Vje8N3bQj+X5G0xZ76KCuiGKUPuxYfoZcGihsocD2jEuAGE5pHHo4hzuM+zMUWV
HYNUJGshu54PJ71l0Z80THdESkGKSQavpHEVcuiSvPXOuMiKptrRfuikKmIc+M7fWjNtfcQ8QiDC
OBqNmoyIG1ufCmh7hmmTZCerXaU0RKhkQytkLsWUPkY0OsgdCzGAJjIIefQrqkFTB1m6dX32AxSh
o2HT4Mk5tViZDxW4eJWktwdFi0Yz3H/WYTcCT7tvCG57TergQ25nGtKKblCI/Exw56i2AL0mrSm5
PGAPeGJZY5fUK+TL/3uuSUXSnBUtCzFr+z6YWtEvwz2D4J5UA7cz4EoYbwDQ5DeNd3opa1osJtHN
b4E6OFhnkgcpvK/70lMt/TspMcE5zC3jnjo9fCXNnRKas9Xi8R6rIfjk3HiQeW97uD7ZbDYbj0wC
kG9v52BPdCRaV0cMC4kypCrd+hvhS8BtO/jfY0nRHpKCpEAp70XUfAORj5j5M3lV5n94znYdeJwS
js/VnXJvoPu8l1o/1dQmDGGl9ExLu4wO1MLAtfvBkDDSfU7VTQYTZ159X4gJgP30LtTYFA11vMOg
T7XaXfPHp6WfmrpiIfOkoX0gfj1zSrjZP2adL95cVElGyP04/Zkiuo+O2KI/4AQpRtKrR80W7AOP
zSUOLZBz6q7q69Sr9GDOdMz5/AKIQ6BTCOORq61RdJORe81Tso+dhdCS3NgpgBpTSCfqLxhd3xlS
QkBxU3YtpcuAJ20loQelKjBgHczDWugl717r5Leb1amTV8j7qjmafaj7tXR5wyU6CdAobK1PeNcC
Rxo2SbzG0UD6OFzt9p5hj0frq4sb+KuzDbijPt3DpqxrklW+H/zvcm7S2166Fs/RJs0Hft30r3R9
yvGbU7G/yoI41x/7VdSrDgQsU2bQABdooGB4FPaduidDE2shy17exZ2BXw+t+RdamRPPIaJE74Vu
MQdDQRclmHvlMOZghGvsI5YEcYQU0mi1yEOMWDEMxT/HX4GIlWLA/uEYXanuwmkyVMXG5/bJ1jgz
CK2im5mIQ28kuGNdIgZ1eQ23K1FvDxso2LIrU/aBFd1l/3qaP07uB+vwHC8g1Oqh0AzFa8Tg+04P
MrhmTe78xgpRxi4qWZ1Nlf5aCdYg+jCsV3ohDQ/C3bY2DnC5wjKPN3+qV7ijBEHp+YQqVaOIt51B
tnCbRwgMlCiuR/2NqXJCQ0DlZhcDaBTNZv36cxWVjH7+dzb9bCKc0nWCyIx1M8xgIQoHsUfFqqYN
55jL48Dkhbo0HU8ZpK8akcFraB15Fsg33oYfnT1T1I/P6I9fWzliY+OejD5+FAGvzn/oBRs1Toa0
JJoqSaDm/XNCY/mjPjdK5geJ4B0t6WzAIbVeSRDVlZBPOfoSyq6A+E5e5jqPiZxnSNEjnHO/ZQ8g
OOZZa0gRCjJKUfuP2914Yfqb4ypgjcxKVe0h9Mv0D3FmLKl8vqgLnlGXDEQu7/q4jvgrJ1puriWk
1SDDxSc3ZHCit3mrL/9prSvsLpYNBog63Kzi9wBWO+h5OInmjFvShKrXEovP4bH7IqhrX6IrbG/c
kCAiRDIha5isVmCl34sVz58MG447YsPYJlXb1JH2y8BNqiWiWAtG3no5qJod3J6EX+FbB9xfEPEC
BIUAJdzUaby9DxUkV+Ua9yIHnv0CS3PJdQkWHd2RkZroU8aKsHYpRKEv9a5ZFrL+zah3NluFQzVq
P/Uum0t+w/MGnCA1JyQBM4rtRw0nkLXOoxjUG2w6MBE1Y6iauRiEPcJYZan/F6pi8w0+wVpMs51J
riv9P+mAuV0K8B13zOLpmEHpndSnCm5By17ltonzmVI00nyFJpOFRESyrHWDUuX6ytfg4XWyOeZD
kZxZ628625UcCitVu6ba1rYlsOzyzOsYPi4O388i5rtBKxK1i4a3HroGyxOV7SSKHLd6NE2kdGAw
FShzqb/PkaTO9f9cK+37PnlScW/taRzl6g279EqPnWECkmUQ4+V+rNsSoL+xRei+d8JEoc8G4eSv
yRCwntdtA2uQDM6wPXUtXD4FzUVNezvfEgYjqZSHtSJrKgqqgEInfReQh8alIcDxD9xr7cMdLrFx
NkyEC0duSlKyMV6KxSovlaspJFOsMlaUwGn7g/UPK3NdSBRfXOKzfgzup0JlO1rKlNcpFN4kRK2b
iDmtARppj8qsIJ44UWaxnd2qrkCmfsJZNupbvYn4ja+5P5wipisDgokYcLkb2onFh8dPlsc7RalP
pwbAcYdAXRdb5oLRc5//kBWvMzXYMu6NSKsRqSGhLldEhWG2lNIXhqz7caK04dJ28xuvAIfw5Hdq
mOCLNOQOXG7HWgxha/rqQUxknl6pUOtLVfnksVitdQyEO3T7XuMNpOIzEG3huOrBwpcg6/5yuQBb
wHMRCsfPj7pXKVU10x9VbOJ9vGtTpikLphWiCVC9Fxa3GzTneGBpOylq2OBWoFhWHUlTGXkt5K5h
PU3WHfrvIbLMvc5kZ0SQHnptKgfIxXL9jyXttl5j1uirOq0I19Btm+3CsoplEw8ak38FEe2mAs0x
HevY7COD69fX1GbYR1hWa7hrwuN1SoZrWtWtuBCIZges17dofLKcLDF6ouOf3Izo9ka4XsV+mv7S
k/wqrmw1ZpQ7n8AqHZfsggq4RSPnqGxuxMHd7sKq1gq85Lw0Ilit9yLUo+YqfpMNB/jpGsauZ600
gaaEl5gcC0cVxisHi66nB/1oodoEymqDf9JhBPPP8kvZwNTOSM3cxBKgaqjGWOi0NmZjOCLE6tKq
hGcK5P1CaJPyN1VXM8G/vOMu9LLmazMaEzytr4L1kcror+6MCFBpSfnWAx74/l/fmYLe3IgSCqxv
ogZsO3VKiBR6Oa1PnylLD1cxNIJ9zy4bgx50lirpVT+0CEg1CfJLpvofyxwVjkPaY9Epj6XJudD5
yLitUcyuihibceOAYypqhJywQPXaM9zu3+J9NMc3KMRyzW/6k4F2QNFZRxezWybdekeJpZZ0Xngc
1RrSf2ByKfuEK5vg3NcLxyIWzlP5iOQesh0fds7C/c21kXMizj3O+8DPpWqvy+kvFyxKVY7rsIhI
YjjBs3y318ho5VX5wMVTTeTVhPk7mnLaR6T3/+u8kSrPik7G2xZ26HFh0kbTvJ/0f+RZ/X830BWJ
9/n16EgJyExv1maf5umbEuZzDmJGFWuvvwW54ejArXnJeihs97bOroMMc4jY+WMTYnBedhUT3zpl
P12XSJ+4P3gEAGZZejx+3FmA7IJFmTgO4/boaKARSqDp8ZCxEfbKAuUCjDb71N1ZbRHUVWhYuM2E
sLFSNGUwVjxwZNQxtj8gh7ivODPK33jcdQI4BPn9Yv+VmRGP395l9BXTm6j5bwBG8VjtZXTdzc2V
vAJVl2C00me0+7p52RN35LPNC9O4AoyYBB3JtzByHFsZ3TPD7DmHGuPM5CEOneBej7xKrxIcHbnc
GQV2ro9TTouOZpdzZy52kLc3urfe4fGUD5p6WEl0mMakhM9RSKNJbz3cGzeVegrVjhyHuEvULmh3
p7vgexQWIa9UcOLpH0TouMwyyEIbLyB+6WjlehWeWP82RXPUFUeXSp6A/dXflmtDb6PbDW5kLpoF
AoUUT5+a46abR2kc/n+3WXA2gT7uOtGcGYbJUlTh2Mi9Ow60ogH5Hb2c6kZOR0g/ns7JtHyk+PWp
CXKbX+2bxt6LjGccHiDVSzsGYIxLVf5Dop36LvlaGHp3MlVrgLohTpQuVFXsBkfT+ad24P+QGBRN
LaVd7X84nBA0iix6FWVLSPczfJlABWLprYKxYoiucQC1YpTHNe083jpoqS7oT2CMkDZz69TrjVOb
v4YP0WNo5VWtrU9TfWWSEhHHoD+F/TGJ9AbSJFrDHWqdNAktY4ewJY6sj1aP1HLOICmcpAd4jU6T
ydmazZUtev+V+pE3+MZ8HmH799hPjHnTz9vGd4XiVoVvhqnuh7wGwk/V69CDSa7/0iK8EsS+kodr
s5sD/P7M/2+NyCLwxsFEG8m3cSSAIjNTkGE2CGdk0FCoQtHFpGbB3m4Fw+IxVBgQdWsODop62ypx
dgHDqZYmDmsd6XzxOSCMEFW+1viDSfmhLFc1iXqXyJJFpoFFPYDhOGHJGkKDy3TnJEveBykI9otx
coSEdNmoX1WGwtbZtkccrvh6ebD14kWfSP6OBBpM/2K4S3qww2YNiEt/BeR3w2vzaE05fiXJC6Kl
+Sdn7PBUIRXMI1TRIY5yclACip9LFszQap1a9DvF5QAy8L8hIWl2Y2zz2oLf0pZFFJhnYhC610UE
e+ZLxxbYiE0KtaduK20f2/4RujhewIZx2IK0F+m3FIX7H4Ep/rosp6Q2Ca1E5Awrrw5jknU3pQ1q
8CtwPeG0Gg7KkWqfdEPVizWaE8EBxzq8XtWyM3q6oi28tqZdQnipoYX4ypMEEv1DlCMLZ7KjKfxM
j1wmdGXXebSYm1yEx4jEUbS23vKes0j/lXM3jPJjymq7f69oLdKX4/q2G+lbe5Jt08RVO/SySUtd
PdB6CMQ6knIGXFveZjh3cPXRSfGRbTkxZxbdows/wE29P5G6tvob7uYrLqrRTm2cGIdAHIgnhp7v
F2lSTRId/9mzcIh93bSosASMFsjXM8cKTWYgggeCNnT7HvSZg+skFPBudhSKowE+y1lC3RvCT0OD
lS+quQKBouyaTDPYNJWpzRqTDS/FX/9bTsPBylHU/Kf9Msl5KMoL5HOWZYPngm33wpQUnxV8IgaY
HoyRRQIR0eg6voFuquzLm96UjCmg4wDawlg81uJbEAM7TbZkEncuCKb5yW95jMGs9/wQeTFuvGtR
qCwS3DXRjA23tgw3MwByW+Z3m/h+ZFRMwASn0sQtgSrMwvzYaANXTeAsdOJCOCrKQNLINptnZsCK
lxnQhIdd8qZTZpGCzH5nMkS5+8PjFxlhSWWkRHtVw+y2TQL/hLyfQi54dviGHsb7xMyof2n6ZpTz
tXPIa16HuUnp3ugBhLrP78s0v3iIz57AFFLFlkGdWjNk2lFvlszNQLhYDo9163DP33fSZaYvcwFG
RjwJeqJHEqFfBkYUAcHHkWkcg1jTakHjg+NqM40lY2TrAVYifyICkUZbCKy/iw2LxDIKEhyZymGR
kqOOR7gq6vF+tDl9WNProVirr2J4/MhFvOCasft8qUpMx3MtUMJitqIgtS2I8P/rxyQQMFCUN6ip
AounftXN+w3x8OZmv1XCBSqNI2HJzT1SGeil7XdGn7vu0pqTWvxGQ2KFYJADIhUXq8IymiC5TNLv
dksb5j/jYJwgzZXZAABPlN6/B9mQ5M/Cb7MdAEAaBB0ZqTdg8EI8qOuLrss0ZOdXfavH94X334dT
IFM3NlRg92c2bFhEQiIG+CZdYbPyd6scEyj9geOsLP1hTlnSwvQxJ0XKdeq1UEjlf/J0jpuCm2hz
MyzhHfqYO9hHpBIgua0CXogArZq7ui44N3sRvbpwxcVLLrk3Df+13i4QihQtVFut4Gp6vh8CbmCB
8UWcG9TNdfQJiMPn50qZ4pc1dfm1AqksT370Qi68MVQ5T8FgA+Sj2qjy/UIjy8sj3B7JMgk/zUl1
CNAwtpWyA9/8tudyB4kpO7bPBJNw0TbH3ahZa7eW7lKbKua74jg+zhV0bdJW1Gmen7ggjIWHYmUk
gAdmaoP8spt8m5ZgtWH18e/+qU/sIslrkR6Y3o+Fs9cba7gitiw7hDM6yk4pPzQIscbo2KSgIJVO
0gUMFt+vdNQwfiVwxCYIT42pfcu3lLa0gltMiS/gpy4EJqrGZ3gNljBs0EgTaa1afp6CDanKd20q
HQGjYVZfhX9YQOdpz+4jjSbg/Z0qDuiAeCx4H0MVq0+RtgXRYe5hlCj5w8YaBHVj4soyVN6viTEi
5VDbHtoYoSOuQFyYhO6VIj+/j2LCdBQbbut/zOEBpDp51oBAdqeHucnFHwjVZNZzXn6QhRTzkpol
6ebE+BRRTrFlYUWMwaXNCi4cd8QiSpYnGNboFrrEmhFJXLqDrnNLYI9QbVIadWC/VXSa0MB9Hp0J
TmhlYkCQsZpZuQf7YfPYWRV+XQ5T8Z6/9ZXfcCX2QhybiecnF6xjk2SHqx6X+Goa5YqlPhv8q5wu
1pYJ2PKZoRnVKNjHxWovjc1ZbaWOQQNsHazM8GC3gfLEvESTvuL/Ofy1WZz+LONSuPnvrvxJDOoB
ItwyxuJALUi90KNILggvKUQZX14sni/OuhIg6T9cBPgdVYBTr9ALDwR9Uxu6Q/4cZXp4M8omYJ3g
lhV9Ugq5SPMmFN7ME2txr1aybU3wWizS7a4ioN/9uWPE9rXdmEpsJuToXD5XnHNVbagkboKkqBTB
6VrB7FSxeW/QG3htFwbcNl3CalA/VaecH3jiMzDiOfvUpF4KzQ0ZeqQKHtx8nEm4ca60Lq3dX7v5
gcfm14/LomwXTsYokAeEouaiPir+FHA/4aqN3ziJ7If7VE6buAbJGvVIBMARlT59UOG+uzueCvcB
GY1zfQiPRR4MX3Ch2bHCp0Bkz0eEg5rad2EydmilnNTGWqtMBrA2T3wQZnYlEsGIZYZPmWimaTdB
6TZGmbGbLOXohuZDJaPEisK5t5LLROyZvC/J3BFVnewQTmc6mHlLUC7vUkrBxxM3fT1OUuDd7TOL
4R5o8YKnc29d46ycr1wBk6V3VEy3g/W499mK0iHd4HChIMJ7m64rXQC5dDFH+fP5d9CpuXTuNn+l
5BB77CqshF8EbCXiZDlNFt1qxpeLSjrsJIE8sP5NTwduote4IJIRHRJSlr3EQjFEkiQ1+DmYTYak
BIhn1/UZbvskSBj4OiAiKFt8vezA3EB09AwwAfiql5hLzvQPCBKVLB131n5XAqfJvDVsNeXKdMAj
2TtpKT7Z03/OsXh+H36oa9MO9uW6fkMq02WydYGgB9vjpCDrK9cB2OSqhnsigVykZypzbNRySARu
rbxnxO5oJiM6h2jErqaDNLxLeO4ZvPuTJzUoRibbBVwZCqnuOibB5SWA9SdQDltMpqDKTiDiirB2
9RiWzPDeEh1OL9ZRclIIh96OIbe8nyBGs/e/L3+zvbzkSopGbjNdgIYJR0VW5VVTJetTRAk9fcOZ
LJi6M++ZrihlECinTg8YmEsdE0GLQ0i9RVS47dOOgnCxYeQ6ZapS/9IUZWAg4BVkEKaFlO2XhYdl
uqvXZVNM2m16q2qp67HDJlV0wyDXrpgrMW4WvSq35wN2Mr7b3b9YwZUWcCty9AiA0BUYpeCzeGq5
i/4UwunwsoZDLgCcmR9NB1/KXtbsSsGaRvH0y62Ak2FEs5iMee7kGQBbuLbVjB086Pz9liGvuj6X
MycZpkqTDIk3St2ftAAvmkg1Ns6C9BNndLqnzoJ+Wcls3/Wo6d8eYAV1epwFJOimdGZGJXYWNFCI
J00qKpn0xfLsNLJHijuNN5ghcbLiXRfwg+z8iJgM3iUfFdGXo2VilxiKjBIlrt+VCtjDlgmmpKsv
Un25213XK/KNAvNPwa9HJpnfBU763WvatMaYvaJeMs6fLZpD4a7FD3916C1nMXPg9n7NfgkyVL3D
+Cl712iGApS9jyG/i1jO6d2FcAnGFBMxeVBS0raWIDotCb6LgdyUMP1Adf6Jf3bfgSsR8RjxgALA
ob9LlQ7wHrR+y1CSH0zPBanSOu8vRWq+vBtNhjZ4Q2HI6gqNhgs+K749+ksb/F2/5NPN5wlNgWm1
ezC2iyU3trkOCIo7fMgXAqu/PKE2dAz27wHZMd8PJDAv6GP0K5AaL3CpKFV1qVdpF6MIt1JgPNcr
kbokngUOYLAoSmRWbRMwxBT4JA+nRIQkJVhS8htq0rj9kwnJZPvvUip84yxtMnq1yW5LUYNbhywc
ghaMVyoVo9gZgff1nyO/JtKl1sC7pTio4vnym2hKE0q0L/JjLWMVnymYJmwUo0vLWxaKx4URCz29
odyghJAPhPa4W0CXg+x3YnzpGWsgDoWPxJvujDeK8Wl7XYEUfFaY1mR6m00ZkgDJn+ILFSLVbASh
G7Zt7MEXguPg/X391eXubqlJDIFzowkfug3FIigdXCEOoHZQFBumH30f0PhFydiht1gAJs+mx9gl
e9rbu+E/yaAS8LCv6KsfzYgyG1iISSZjGGG7Uu9d2UZ1DPwicG7ivaQqyghGrzaJMbkBpeXXufSA
CU45DP+D0LtJwVvAOe3r9xvuTid6UeKB7MVu1PyAAcD8DHTOWyfo8nxy9ndS+UTVh/hCTaslYpqt
tdRfyBCKfIpFI0KJMyOhIk4Y0SVfiOZNQax2VSr7Lm7FPSJGUU+2rUHrfIZCjw1NesAmrw7wNlCn
LqC7rCoCiuGfwCDLbvlZ5XqGjg4u0ZK6Wae1W/jwd3Mnqrq8kdHdZ+iMcAkLVUumCw9HGoVp6bC3
b43sQc58USgTmanMyODWDgSRg5BEs3DE0PEtMDJgXry0jQp4O3LGmQS0670Nnp6yEXtWeMqXFMqF
X9G8UnPBK8tqcLG01BOjFMohaX0KD4UZUwMnE2imnDgAdIW0Ke3U6pmyRHlXFEeCviuI4j/tulf0
idk1h2YkAunv0WNUQSk+mbZJvS3nI3Wy8PhJBRWX9dl/dV51IQzAzWKFpt1I+nb2+f2gUUv71gda
83vYVju4AU1pUL8DqGmMUjbz3y74VEiuL1o/qX1p8LQaFzfA8+Uji76LBiRQkhnZRxDBsc3cjV6x
w2OwkjlVz5BjS2A7P1yske6G/6MZTBXNM2NgVIvG5gAIbCDcxwasmPyl/HJbAZHyhbGG2kjihCBm
ZHYxZYuTQWUgCljFwvl2ZDEZiD+eQl8XgnixkzqY3mc8WPDg6cSlRbZym+zpnvKm5idiPbrkPzd4
ECsRYxfkFOMYeARCce32o7FEMYhD9kuJcyxV2OuKd1DoZ1mUVKsKJq5rFDMOEvhFiFi0kXj0xUCc
Ueh+8myA+GSDivOZkgekehaAqE6vFRr+R78H3flpNkVxUuS+lHnkG3ZHOdV/r3ihJZwt8tHrCIx6
gAH/Ug/uyoguho9sKRKmaLSLTPzvVCtyuHkc2VzupWED/VPil6HtCI1qXY54vcBa9v8SpAKuhfat
aWKVbqoL5HEz1GhLGaOauZ2lP/qzUbcfH1pyDfIYgRCw6DTAfKCWiRIfVPcyi83+F85CI1xsfQhy
SLapUja4673aqZGYpNHMZRERjSZ4lP0ubD78UObrzNw0ZoDXaV+SUdkSVr/2UhKOSbTH4WyZfInH
Qpfqc15NXNW/f7hqfDnaRQsX+lm42RJngKKGtqLVrw1iy7ErF/6Zq90b/8cnC9Uhmqmh0U9IYWaj
KKsBHpbAvf3naWLq1rXyWu6Lv5uuFXhPmUS0jTdIZLQcLT52sOS7o0yGbwG0pecKAHMEsfGvhdRs
vJJjk9l4RCqoUuyC+QXrSyqW3WrVwknDWS3gPS84JH0U6gDdum6JLedrGifeyU/u9W8K9L2dCNf8
UHjPkIdRLIR/0KILk9jg+NsiO7rgfE7YQ9BpQ7i8ik466UtYNjUIDY1/yeNRrxNNV9v7dLB20OtW
zyIXgZl9qku6aCKHoZafYxX8WGdMhMCVuuX6nrPh1Ptv85qjc2PuwIzRE7REVg5SP2vBD8Sh6IwC
0yhuOkFpbwxtZuXDgOnOhDJPJjWl0TnyaGAawBnSnjGckPLWN3qLAKQnP25IA2Gh3guAZFBEXdyN
LpabmKviIsZTzm3ahUmebBXW5x983nvS4tCIibKrFsoAR5qxnIcNKmbFm+ZmjsRcMJlec/OmYZzl
4kEl9WqN2lZuIr//QG4qd5OH3AGE10tVwjgHmYF7y+mPkvOSuRZSGK8AqBydpw8p9B3LOXgMaQ8a
hlrG50V5INK1t59s5cvk0ds5dZniC6m4Ju5z5THg8OkNz+5vLQSEeFs0lhi+5CMrhn0//63azHv7
a9i7/k/VmiwRsOQJ1uFfMJpP4gkZsnPodPgxGIJDK55Nv1d1IEkHbUJ5fudPCEHkc/SsN9CLnB0o
tyX+Wgv25l7DM6jqje2QEsTl807Q9uT9Nndg8WzNKZmUWIwwp8uXmG5E9RW1g7jyAvwUcfUOfacX
OHuyYZlcgsc9DdODPCV+bgwRQiBSZS4EzPN0n3hGzFDLav32g44s3tsD9AbayWbfMtVo4LE170pj
oJb0y1ExEAtrBbfO2JRM2pjJWq2YFT1FuLQ9GtSzfc9izyNKoM8K4/og0ENqFKaelO+in3zQorAn
Heo992xkgYP55Wp1i485pBpAZaTUoz1OJroSleBt5R4xNh6LEgUPcajGssNvVONhNz9ZFxJmRLiG
cVdApZvOedKrp2DSMEIvp1lAS2c86FkLKV/UwVlx/kTGYUxNScO+WXqkdrriJcvuWE6iq4SX7FpV
uVQe8X8D94MLeCbfG8aX1+D7K5rEosYyO9LNuM3mS87j1TRVy0r1k5acVGhEN6qbOZaPlustuvmB
qyXCSLE0kdGrAGMBH5pSymegOborHty/Flbo/6+NH2cDLARFr64pX8Zf++tzmMyMX8m4PCL9nq76
7feVmacfEHDfG6bDpoKODjr1o7ksd0Heuap9iL8qx9pX6yIuzCkrFT5ChA8M2wBsSdGyI6xInNPv
9zH15xNS72E/MiVRoZBefRgv6Q2U3rj9FopwRNvFyaP5buZXZAYHKaPkQMSjOMVbvGE96UHNc0fi
VI6jQyn03zf7eGweUF8vAun+6BklH7zg6FR3BIko1UF0bejcVqD+Jos4FglDTs0L9QD7sCtWp7R0
RWTJ/2v9jHRyigCAe/lb13DNEhVKIPnswmfGCgYpGWbF+aXpAL8HjnUHNCGTIY8CYc5pDBhZIIpp
ID+LqPisBnavBg6hgxF5yxH5HCwcz9PmLc1lxsv0pQLHge80bVj0wVGHqkKbX6BAJQ/BlEmI0ClB
wJO5mf8u81rCXx4QBzK38oF13N//gX/vPqz2QlvdR3DPq/R5+8bnU46qsYmRe7c/09/JM/jJPcUZ
D9p0tecZGbI8UHIhvQAW8i5IETOxUF8DoySmBC9nS/KpIbNkpE4c8McHZcIDPxW4PpdnvXVqPEvp
oxhRKfvn9hDwvgAIDpqNf84laFlnb2LMBis4opVAhSepm35Blvi9LVkAIxXwYUqs0dvBwglM8P/w
MHItw2LkAyYTnaZUZrdBg5CZY/Df3nwEYngHlSM1FaVaCYDjESQEkK1rY5auN/wfHKUqG+WWPbHc
ksK4tiY1T7bNhki3FQ7YqGQiPVQEIgDi2Rd7w90QMom3Pr4Abc9RmmYycKfLtNlJ9hxLs4SBbWR4
oueDC3ETxh5U4LL47QhDY5MSCzWAnE68YP2OlIuygnGsHV0onbjNAPWoyEP1J/DqDoXiKbYBBDBQ
S+XUh5IpFlJ1Wh/rqWGZeooQQ3H/ShawfNcPiGaVKTjyb0+Zm3eWPEUhGCWLmawAbC4g4auD4Cud
SoYLMw2rjvCpAgR+l3FhpTeZXiZ6zeEfCW0RrkiZesU4jVTRPl+AzTiJ0Cr+OhNyO/ajfOGnZNWc
A9YMNn8ntIo0/wgA2SVGOdVcU53ill9dAr2K/I8umgfG5oyZ6WuDaJK+dYacDt7RZiBcJM6nMRio
Z9fTWzrDxEifpq8aeATA2TM0K1Cg/gU8LV9CyBwDi0sYgG1PG3jpRMQZAE9JF0we1MVnupk7T5m7
SfZDDHL4AWmBPcn1va+/b8mU6gwbK+XUEXD1lKePMDE0nXBoVjjYzLws07y5WpPeaQyK9UUXqh43
DFXaCkZmzN86nBDtAndn1bqR6vrU5W2acapMsX+1TE2rZm+LkH6B00381qXo8HtOmzRy5l1arLZ7
kp89A1TwcMJdWFV5CjNYB+pnCfk0XNrJmB/VASOx/GtaR+mYA2LoZ81dprqeJHN92E2KXDD1Qkky
AIb5gQgAUp2NAnZBo+043ggRa4+gc18r+CRmXtR48CeF2hqe7z7fbFnZ4DpKFRYoyIhw28ITl8n6
KMqnR34jlDKLR19dfW+VEZPR9RSSDwsCSiyqrVP8lqBVH8RHQBpxJ6CiOgc1XyNKQ66uu/m+zLTO
EaG1VhJ/geuzYczsOZxz1bwd9DKBtdOU/GpPUcGl9BHu7OXH7BG5/ULBXbemPIHJuVVbQmYsMpRf
qrvExuf8qH4LPAeWzasMxRhMUSlKfxrqOk/9LkhOkE+XgMwXyxuY6vMwQ+J3YF1hDmRtjY5e/yHy
FfJOelhYRlPQAQ2mowQu15CuHm8zztidSXYwF+/YvfjZCAgrqI+qiV8P72nWBJdh5rnBzr40rJBS
bAF7whlPsFhXRD41p+CC8nt0ghlK7HnI9Vl73XiVASZpukhFmpMkS7FXHyoSVmvnj7xp/Jr3F5Xe
EgH9vRZHnRKg3Kz0BnnMI27SB8la+0phqn0v1Z7TRUOKtYZELM32hkytMi+B0x7+rtW7a27YfBrf
LyEFeAedPXWZ/SQ7DwX2Ug/Nx20S1s8a4eu2RXkYsdgrpExI5i2N0KjED96eQl5DE0VofeDQhqx/
N67kdF0MdLRC0I0plFqnnSTTKCDdAXo/53j6RHaNPrc8l2eEWChUNxiJTmAF9NxYR6u5TXMbTJHh
YURz2ZoSPBeZ92oAwG7et7i/YDrKWQQgpuq7EwhD5jiVQfsXwrS6JZsPRK96rnzu3nroldB8jxur
eIif9ScGBP8EtDlzcthQnGvnrxxtXAXhY985OExYRFuIAtZg5nvQpwahDSyKchtbriT36xYrTjxo
Ul+phQR/00cfFKEZvfltOJxPnk/M34qqy14Kzjx3glO0XisKS7wgYrtvhE7y0iVFL6iM9nc3fIpE
8/rSwYF7150A5PWqKGLsXIPZgXceT509xCsy3hXs659muZoadv+PyOuA2fy7l6WctLLPdPmYUEsG
z8uMRwDv0vHZGAAhfbx0puyZee5Rr16ZNhOWoJkvISdD+3uSPUWsK/yDm9GqcJPfHz02ygFN9xI0
fNansJ5xjBgYb/WsQ3Pb4+GrTQk1+z6fu2fivdg0TfEKmo7nR/RG0iE8KdGqw61aelNkDfKpoIaP
L4RgzVbLGX+2R4lFvbKi3RSGGV4qooEYAOErVkNmK5QOjPaj5oOr37ucRewezS+LnXbo/7PF9ExJ
FGb/3QyHNye/2KrkTR5gwJTHDCkSHBbIU8IArS4iuZbdtMPWyyVQSP6XRDv3JWxO4gMj/T5gB4SH
4DRTOpz11FSAlZkHgKIBs2flIkEz3RhHIvVNdsCxF8UQss0OH/U7xaxsKQJefgeCKt+O/bLLWSOf
N6juk4G0nViEoUaRqqp3u88kXK3+qYm11kPHCGtoz+xipFVcWA+FxI8mO4pcS9+tAVU+K1oAy8AB
gczHe9yyiEgk76BGcoANcdc954JWbfZVcIBa+8tIjBUL84ZG9JOfRlLEGMpfaUDuyOwyDc1vg1gK
CEhQuCvFN/uWyB1lMqEdGwwx+gaTtI9RkL7d8GnVlxw5W49X2TgxYOOmYEGOYkY4tMsJQyTNpFZe
b+m3irE5H2I7Sja3OjoYvCEj/JnH73O+yw/utOIbvANuRBt0ZJWaKCDZ9RihAZrj7JjCvFP76PEg
GG2R6Hsr1Fx3e9afjMQtqW98C1x954rSUzwwy0JdUl93Eg3II5nn3RJBaI0sOpSUsaX1LoqEDXED
YY0iNCL3CQDgxA7wh40SByN545//7e36WVRWzHMydFbPYum7QA8PwaxevzeQoa3g5MN/uZzDNpS/
uWhozGITM87Q1WzuQCv1vFMDeEFHuBkemYUS84BqX8gVPVyoxKJTXuQ+XfIevJoPJLopAkZIU4Es
EC+uro5HHbHbVx0zsOAP5qw0ajYXUIRjB8/N7vf+i6q2I9ODQH4exPu5z0M1Kf4Z8gcjItxhdGcz
ov7bP7XxrxJZrFRo8Zvxy70eCyFF5a0aQtJxDinVl8e57DtwJmWno6wGOunu8M7l2TebVjuQuzQP
0qSydfoikhSP59tDBT9f+wdXnHuxOamXhz8xpBMhDs8CKMo9s+s+S35RNaN0SeRSwnNkyrbBgwTP
DyC6FnQKQJBEhTIUg3OrxRR6HNvgkMXpRsHPI8UXkgkyPsw9N3Vxlf0Bd2gHLOGmHTzYnKj2jOvi
fsEQLhkrPt4RNLJEChhustdJNmMoTEdqzMif8RL+Uniol3m1lAXgbPMK/OH1/EN2lZnNobLBg4ls
yZLpKqU6/0II5/788ARuc1/6Ya7yL7Zp30NspoT9ixL+2XTmKwHk4zltHXFfmspVotxYmzKdnah5
4ypJ24UEHKoCx52tYMi9hYVqnbpSTuJPW7ZIA5bpCpTbySt/1GbEEkwiqY3IbuQjP625b+o7LelV
72YMCt2hDOcAWx+RsKUTQ4c21sV1Mh+QsE93O6BMMC2/8mL7dQDDvo9N4Vh0jcWXw/0n5sT4FLxB
EeO+VXiKAg5mkL0wqXJgVEphlkNees9W2Fe4f8yjnRK4PYjswI83R7dT6n7G/45MT/bihnAFmxm5
ZXGCvPkBJVzdtiMdEOTUtzOin6qCKdbVDXc6kSLjO99/cEeRvCCkqxUXLqh2VaYv0XJqPU48mGj8
rAgJXXtXbyaB5rPIQ7X8zgBMHZKgGVTHBZMkIWO3wuQML3qMhKWqXtZp0bsEumVFBAiEJusFFEQn
M4CAaBkjb3X5pEyTCqO1Lxs1t+jbwfcddsMdc1dJWjRqw8H9PAPEjUFnsqFvL0hTzC15QQsk/DHT
bfbpXljOY0mGELHZticuHGxOXxwJMnXc817f8Gu61x166IZr2bJ+0KHBas78tQ7gzAdyQ8ryjbDe
M304atvxAdO+pN7CZ0nkREYsToz3fl0Lwj2sF/d7hOAUuApkWj7MnzqquyvNiMO0LJJR+kxBjFAi
Mq+kZbPI+TgLgsWxzvHpaOOf0kTQ5mhlzs1Q2s/ZRIROr09XpwOtN9ebqD+dQdnJPQuRQsqahHEJ
vUAOXOUmmBxQVCG3CeCZyrkQGOoy/SXj/Y3HwsQAHMGwkkE2ElRbdcLVb9zg/5qnSsMGoeTEDtS3
9xVGD4w3qSXib/pfjWYWA+Z9mJpySeKDUi0Cd8ydbsqIRjh0rKrwVzWwqZkPAu6nYJKjS6QS7/WF
CytyMKDGYqmUwDSJw+zVMufsSSN0iSdHdDNUKrQGT/9adxKJiKLhxOYbAC3zlFT1Tct9xOy37BHc
F52o6wDfUaJoBWUSHX+4rLYfmiUYtpr+yoBIC/mlhO1Sjq3gkwa29DpCD716nyGhiyhGerQ7VOSI
Hx17hwyHdzZA7OtvnW2GpGuoSVsGWtzQWagcz3rxsFn6RkG+w60bL7swdV/z1n+XPhRNlMS2brEy
sYLaCnYVItY9AF6Os/4j/okTT8J99/UK54M6LhwgPlxZiy7rScsBntG3dv48tPFtgp3UlkuLAIXV
XetPXvKHmJtdHG2oGRLhzXr1idFsX88yaNZu77dD9Z/08PbhxwDlLSeUErBkXAUspuSiNXMV1iKf
1tJ6ONY/H2EU8bHQjzjagORAo+cJ636Q7S+U7E2lf908D5gPQ/X3CWPzw3MuPX0YLuWAI9/v7EgW
W1wc+xECnnJEVcUJA9jacywqlGdiyrvr9SO5TlOxsWCFojVs2LlgLSbFcx4+SbcqC6n8C29FxLMi
FYq4ropQ8tnRaf8dMKT0BWzdDO/wIxGuSGaRyME7q2fy3CZs1RKMTeWmkgm/PzsFntzCZS6+8CV7
qYMFhNk1udNfX9vh7zmWRLdeDVkprAvVlgtvedn3xs4VOrejxx6EPgDazxeZDS2pPY8Ucc3c8tPe
lONGisyp//6mxJeff/VTaQNNAxyWC3lWm/n+gmOoDEidGjQef9SPaxvs9NSMNKGDYThfE0Vhxc/6
fXXBmTFpoVy8TGEyLcU+/jKScFDU/p/DqKCOem4qRpclG/19Af/JGo5K7uKYsyHMJ7dyqI9xvD4A
fTlz2R/dTvQWEKjd8SE5ctepMM38Spm5vqL8Ng7zD8pRa0n24jD0t/fAVs2y2fLeW1LizbptTSW2
7Rwho1qbV6VF42FVJZF/3lRDSQMpsTQJcPrgsjyi+jTrBbMh+mhfTutH7B8+a1ulewxZHlVRN4Rh
59+QS8oy+2psTXm8UOZpnutDm+r952HMOKKonDFdW1m7oNfeb/dmKCIOWuhsA4gubNRg9tbViy/m
mT4RqZKUdJDbSA5H0+7yjm/ateSvspt8LMLFBYConARJsgcWz04YK3SFdLplPEI7yWWGEc+Cu1Om
8iIFF/U/q1TjYPT0TIHMTtCe6uoitgOmRABJdjv86fEDQWskAHLp1iYyQOX90Eg8qp936uUPt3Aq
L/euW7KMq38hlqy6gLNoKMYPZlhRVps1vnT/54mgSpwbcG7KV11JRWX2Ot96xDBvooar+u52WYP7
krqll/R4sWIdiCaCJnTOp+IZGUJaglKwsm7FTygWDJDvT90uH90nbHnvpW6n86Oo/7k/N8AmmPku
vF4oqtpjosiu/3LlOp8GV8dA5VAp4K/3yDFi6sLga0LvQEO0bIYwZuzDiv6pNZPSvm+Me/24JYXO
+an0db9GzviAoI8B+VHigx4H/nC6yRKA7CUhcK2JghFmr7/gH1UbCq9Gic+s/PXjVLYpOCk/szig
j8D4TyaO7AEFTU5+RP9fovzbHhK56D6JB8QIEaWbH+soB1V/AwELDfMmG+P+PQl40QBQaP39+6yW
YzfIAUfy/qEGWu/OTHqZBS5uTL98XBzCElIx+Fc3r7m62SHrOlI2Rl+WByxrW3bKCQhadK9GJTm7
QhBdQx391ybs2C0oFl7H2Q9oJ5Dj051KHMbUP0FAt8qpPlUd1ichMSArNl8Rk7DBT2NT9ecFAV5o
frK3dXnQDMQNemY/f54ewcMhlbg9M1cWELK12rpw9aJXV7K+Y/VtiaQnTymV2vtkWyG70FnrqxwA
eOWG32p/Jv6P5obPUuQsEyNU5zjqkPVFPy7l3A6tEMZVlgg1DPpOu3/Ra83tQCzjcbO+ANsTqDhj
Pz56LrXhXXoqj9rmiWAVwQyu6ypuBOFro9BrAkNljU60zY5lBQR9ErwSTRFL9KHkPBqcVXyIzGPc
j0uB9FhlCLtSuwNRHijWwaGm7HaIzgmsbzJ+HUWgmPWokJh0OIyyml7Jh9FBLmnE3YTtMWivq2g7
wOltTgYSR5iTU/zKMrq07jZt/WnTY2r2iH0xdGuWo27dlXHgBP+EGJ2bgUIx9u5Ujc5Jz7/ppC3y
4jXl1JzB/YXjrPtwd6sC7Z0QQgHgKeefmWwEDXRPV8neS9O4azs2jftufLo9pI4COVrEj1woGhVa
tIZRdC527yC2x673EYve4v3qvqfkjWnGPXj2ZYXvAUrp5Y+WXLy5Nt9idwkmnOGaJzu8g1qNi7c7
Anss2uoD2+VNWbywSaXlNbo94HXuhVPk7W2VJTSO2HAmbvC0J8rYl0qleJIzDvVHrGqp6MiTgbsZ
v76CPPFTYFKS4onkIR3ly2RdEelsLVOyWVEffdRE8qk7htrHidpYHnu3tdgH2nivRxCkcSk8fVY8
Wy2a10K9ac8RIIoAyRxD7JyBhwp53wjKA0Fy5iTjjpNBIIHM+/M6F3PMk+U9TdYp/wAkYN/qPkxH
9hG2HvhZxO7b09qTBc4gJ8Fp/ew4/PRVwp2HLB2JMWKb0xiiU1JgczwFwbJnINjT1+54RN2sPdRA
rWz5N7FnwwyofihZfI1ZOyPfQouHAwqx60CVT1UXSoxA8yHGmZVDtAuxr8jkZVHKNK3v16KNh6ye
eB5Irpth2LT7461KmA7OdrU5JJuEkmIgmPZpAS0Kasqn7jL+5l9CmRwylq7R8aX5SdkU28StPjad
PvJyIPa9gi/xMvs9JuNobL7Ng1Ofzn4yXNOGot0akM/PZvYwtMjmyHDpyueDhse24d85Lezl5DbW
Ftg5Wro1UJIzg+DP3x1mGDvRfuIbeoAcNgAJhAiaC5tg09/gNd7ju1yCcURi21aMrpCmC3wXLVBs
D8hed75lkX2/bjSsl3darj43QBFVA+/QVPQXMffBZixeYFxFbb2dB6qH8Yo7dQjoBp4b9b6P3K1f
QZAybjCpXAgymZ8RPEaDhnHLi2A/RIEk3iN3O1KT5/9RkxmyAsV7U5iFgFAwsLzxO+XPMaM38EXR
swKUHgX8gggtvuI9EE10Fdk/oV0xH8Syk0Lu0ygTWKpEEW06mcyPJPZ34FYndjBnhbhDQfwE+QyJ
m2Am6Lb1bmNIrddgtBoqF5QaXQU+ZuBo9UOtmTpBKvjJIx0f3CnjuquoVg7Xr+V3c3l698n7gu7a
IGXtEoVtxjNUk5poHaYezMbEIN9q4QgvEXOxhFPHqYpSVv2BudHv/4BAicuQ3lOdXJG9uA97LdVi
RPPPIpYBu24tt+j3f9JkrrzGaJHBxH6/bntuyIcHO5btV6C+wvk0DgSzQAQT09m70XaXO7QheT/l
/d+kFJWa1tuJZX4TkriAIUNi41awnv9mZP3Qp2bTvFlpTbiIlMbebXDcITw5qQ5NmofEHFQZYIFn
qMdSDLi3cfYEj6IHTr7FEJXAnSXCxhXMaZmahr+pa8H/QBc4L7Jo48QwFcqL6Hk7QzxVZ9odfcOm
m4tbwjZ+s98SWUh7OUSX7CgtvhanAJIyayXgJlN7tghD3fwEwlivIz2Uqsj2FbAnTO9QrAz2Ba3s
ZhCRUInDKfBKe7rXAea92dKX2zyxtpYcldWK7O9MTRYZibc0ShrouphStfMFQRjk1SyCvCURhwNt
q5WHBEevRrQ0zmj302PtgcpzthMSHiv0ZkpmpcxgrGrR5ROWrcJEAMKlEyOBQYR/iz4KlpDCONa/
BFU4ONvibqj9pqbmQB7scbskWO/UlhVEjflX0IqYR0u2aMQ6voj0u0No5GqrUWiXehMI3J+2T9qA
WBWkLJoMum2bEMnCXmLOy8M1AHUaczhqSQ97zDZwL2dxD2kJ9G3ZnlOtKST/U0Ohv/FEJ5x9yhKK
NFN8CPN5xoOxgyetdYILHGQO1vDM0jthu6OJtPVk5KNFvTKBfcvT2LfpDgGceZRWVT58M19ZtYq2
DCBof3oSvibjOk3McMxT2xAzPMODIksY5o3k+CxmyHjeYc035i5OGZqJem+ntP/Bg9yvPRoYHQJK
+ygUGNEjmX3nVW+2SfNWv/yqzEIrVRjf6JIXuxN4AXPGz1tRPygSCbFal3fjXSGb8+7vn7IgdQOE
ppOl59hM4mrarPuUx3HiBoR2A6bbGqPD7ThrBMcwxjTEBR83kfl0Z9WOFuAGcBD3STYmXEsWEPoV
DY1//2bz7dYHNIGF+WC4OnKj3xgWq+02qOabKA/Rq3CNE62oNYZgwcCFbkEg8WMyTv5HoMVNlEGC
42BbPy790AyCRtAEca/DrNL6ZYyaa98eTmHuLEMTrh68gQtK5TOJ/LPX8X0BtBRbsJorE9MSEAIX
bjZ6AKc7gIY+6MfyAmFdZ7cJQgCzH22xC5X0+V5+H3piQAsb8g+vupxfjolo7qgGIXQebKvca2XF
lmXnq+JGRylMhxSNpwNb3txA3/mwvLK3snuaNthGY4+6reH5gjzFs2wq/Hsl8tVfnBibaJA7TjaG
bIqfyoUMsTJNhvEqoiwV79vZ6KlA+MwBXUhjhIL5hk1kHqE6B40ANKjLHiFJONmTok7/JUO92lwg
HTR8X2eh11NjhNfPUbFfPitRVnj6lUH0em7LehFp4C3RLj4NCvfCKczxzfcxXgoV4pj+RWn65Qm3
evqsxHM/Z2HE09k3iMUFH3YFjAsMXHDNRwSpfk/wg0y+HQcnSSZ+yKPazlVUp7gf7P9XYG2dV35Z
4ZEfslfl0+wTe9c/WNsTIKHGT7cjhXlbajDH8B6k4JG9W+Q1l5Vs1wqATWu2SHyUtsekty9SmBZ+
SEF5V0g4midSFz8hvcDHr7JsDAZaCCp91amAjsCpFXM9XnFUwqcXIzQes2DGH0ypyNFtlRL6RBDr
7oJIt12xdYN89PxGC4YyiwL+PCi7yZVe2OM3ELGyk8o6dHsfCwv3lWkvL3cKcIkDMqC+W3mW0UgN
kupTfslFc9cH9ZtZZ+ziF2j9S6FBRo7trr32x+TVLSyxwuvpTe9szmLjqRbNt9QIv8i++Reu8AtS
ErYEey+zMCWkHeolU1jP9dBXPygDA4xuaVoC26EKxjco+QJuU4Hw3gDeKzxoyKFVCuDeiU7GBhDS
2lo5pV/q13HeO2nVKCx1H8+mcFx1tzxIRkHKQReKQ9DNn1OpAN+DAEnGUCJuXVFFEugOe2U+l5B5
K+KifkvSvTFsXrd82yWl6yoyZcdoIgGnO2v74ha9ElBzfEje6Jo4F8CmPDQyeVV9FsNzW9+70eUU
Fvr/kLDaSKi5K78hIEl0HnK8zXVrSBhBZVg5Coi1Kap4YWlYVgrKwjphlGFLCCyNCqlfmYkiZkDk
1jf08vF2ql1ZmYsK5MCpL3ghF67gJNfA8vJevKstN7px0GUC0+/abuX2ScAzDM96/PaG/d40fGdI
MlDGKLOCsd8j2tN5hnH5vi4TVofQExJvUKlGFM226Zijl4WECnk5knluYzwTIs40k8oyV0x5FpZr
sGgm+W1jEWujRHU04Bq9+1zuMHZFJRRoZYeqA7wSbR4To/XqZTFTHWZgL3OOHh1LkjGgro1EGnOj
cI9ncmmifg8G5T1b94ph3mR+AwB4ohk2/aCFCQG8PjSqCmuEkyCDM0yIjAOXu8QBUckmTF2Xq+RR
an4Kqx/ZIytbQuLvnWxgxT01b9tjLtLLWeDAr+sxxmDURN+yCldhCOOXhm4l9K/Wj5C9R2Q9MGOA
mpNd5gxYt61QiyelTwlqxgirfPMSNMg3nAPIkayxtSsZLoP2WrCtJfdLiiymAQ83swi2UGpBX/XR
JrGHC4yv7Hk8Jnu0lAPf2+jX8OQYNtBcqmEshjykterILArTKjdiBAtSd1S9KE0SOLGRac9Ul231
/cLmds8RkuUWHLsS95EURkwYepCUHsxFpUdTHCEWHSdlRTnJUcqN9cuz6HcslVhSWGEpCdHVGPXy
ubwHnhoCZ8bqP0hXNiCLoWa6jTBxDl5AdXitkg6lF/Sl9AbHhKSfvKf8HYGSo8DZ9NsNh92+X3g0
gFA8FJHXbrWy354qivXfgh5kzUU1bwM6pSNdvk9eJ6Ohspyn59wGla8hXQwF6gB9MjTXEFHKpEOB
6C+vR5ncP+TF7JrtxZiufxKVgwaj3XOQc46aJ7vazI9kRL3EHHnwW0bv9T2bmExw3meksSmTOQGK
T6aPr/16ZajZxePUDp7oi/6h9h5KfmpATYowkBajhzAlWHJgA7EMnYdzkNj/0QhlrQ6erWzKWLuE
Jv7fKfDnV6sDBzF4h8Kd++8iBAjm9INytx2Oe6HMhPb1pXs5EfwhlnRQXUmizbMU1V6yU/TrY1j/
OKTRWIe5VpTy3CYWny/4XDotcAfYzFfIB73LnsNs/NTOAeQRZMLS4XFpPDsOxmZJr2L5yjZLVqn+
K6SJBXqQwBUgbS6nA7Kj8lZEqhGsu3Rl5SHkYe05BB2m2KWB11hbcPtkjQQ2LEwtxmJd37E4rBzC
/Iaf2kX9+WGc9Z547/HmlRO5OwIVpJH6TQnrhQ9SEKcx9PK2BrTWSiWlN0gqoEmA5Zdfar7u/P+2
yHQebASUG61+BtFS7I3Nikc+ggPCUGSFLFThjzwVxMYgMBTCoWimMlDgQPfgst1vPVnYdYssgMcG
hfe5duYIcBYq+5CVob/DhHkh0xiR2hW5qVE1jDuAqTT9l5pXbmh1g2Jrj1z7VPL+W64gVsjqEv6e
2u59p8r8BFxMEneKRO5XxZnU8HK1i+q2q11CgoBNziJ/u/n33GBYEOnBXHUeUIFpCwxV7351a7Kb
s8mjtRcqBmFHRjA7MtZs9pUl1DRIdDgH1dvLbCWC87JylYbSi8/fnAxoeZ1Cn/AWY2gHCChHo6GY
QO2CKdOydXttHZE8dQa2skDRLeCkABW2CrFLZl8pOBM812Zfb5zbfiDf3BOO+7vvbKVlqcHJCbCw
A2fFqVv71A2DE3Rls2DWKn4QUcF9W7ozpK2esgi/e1KMdKs7m728M8hheFVqjZjPoKAWbjfgsd7m
mmLPz8+DEaVF8+PzsWdx1aEkfJXFJrZ7EGZbV/TYLviRyGJqx0Uz8EY2PgioCxp2u3sOc43JgpOG
SVKxT3R86HCxrtmZVNZIuKuhoP2glkYFQoa1LNGS8KQbaTwWeoS4SM52N1M5FJxF3KQQrMJR/AT7
ql8QSG3V0gYV4miKjvxK7JMV4WoPNAM0M//yxERmmy0CvvS9Wa4RLghN7WrBL0WSMy7edjkpaVwT
bfdtMgC2LTgXc+xJJQq+004TyoWRssJkV3RCONofd8nzLG9WNYisnwubBfX2DEuLELjAE7Z0G2oN
fy9Reyb1eZquO6djdF73HqAnfG4WUVd0f/nWoAoQOQS13KEDGWTdzC+ktbdgWjcaVxra2H5CYPM2
DoaL+Iyg0xPEbNeYbgpemiYVa7MHbgDuRbG7SikdGDQCiE74t0tSO2haRhqY5SFDTRD1k/fnjmxT
vEFDfeA3z514TKUFJGKkdeJzH/O/28rdB+X1l9Q1MhcZnW8obGb//lftwUpJF65Z61L9Bl/Kc3/t
uBa+xc85Byy3Svtupp6/Idw/ge1Vx/aTvtdw9gK3P45xIXg1cAvQMVeiFGu3W8qFoZEpz1stAPzb
CpBpnuWlqq1olllP2CSI6pll0FKBrNTdWA16KkvbDsamM1C865kSTdnOvbo87PySM/knjIenpWcd
6VpPEwJpRdMG6CTp/DXSup863jioo0A3XhEygmdJNJ6Q6NGaqEM0wdIBOwNC0ZpJcBHvr1TOhXU9
70GKlmCAmb4xdBODOF8qy3+7DLo+hWJpB7PZQgOKwrZkWQkDRa1OfSheZN9ui2/+sEjOdJpRG4gz
L9vLiLD3MzQuMDHPqkbOkTIwxuIQ1DVRYbHmTVqheTZXyB3Vaph95zDiTr7qSAi17PGj5iC3uJ+p
ueY4NcNdyHO4ilgviHaNFAOpIw5xYM93UzP/K7vrLOYz6YjwrkLYWwIoeDCOWLamQ5O6y9BVe8ZQ
83EYtLRXwf0cElM7ezQ7E2KcKpzhYKlVE4Tz9CIRt1rCE/B/Mvr7OcwZlSI276nVjH7Q3g16zA4r
okmik4XWUR20hqTd9AEpZeoWNTRTZ9SGEUVkN7u7Qr7Pnw1hKxY0Nj6D8WJqeJ7xjm8EF+2FNXSn
oEthiJGsNQTuO/MG+arnnr/+7/4s9pQYLcs4Yh5swfzoTI830T/yRftcZuqLXz1nlVEqbeFf5VJ+
AwBRTMxsSQT7Qy52yT+ktAv9YoyBFCxvjiNhrPS7erYIGm82zWpRH5GfURPrpCUjshbAwSXFzhO2
b5Nh1t3m9s7OioDLBpVdTI1OJngl53VSLb4wf4Bt0fTeT2UNSXl3EjSFDa9zl+F8MdQlvDYg3Q93
sA8oXf/rkS/I4OY9pIKCoAe7chXse86fsTT54Je40nJ4+st7VlYefu+frMgqaOxBqd0K9wdo1D9+
/FoZyjeLw/T3pcLnb8mTVgfHy/K3ZwkTwrEm4Qm/SQm2Fvs/KCtLLIrToqrT+fjbbrjBpTNN8fC2
4wPH7m3lfZzvXkCZq9r+uZSaaLnHtlOOU/hGNjaoleCXIrjeHkm9EMU6PFQVPZnI/hYdVmwU18mG
WuIU+xb8CzbD0wN0nG/OxoANaC2wM4VsySyhxE6SkzPZKAiWtMGsP5pS6/R51POmox5R5cQTt16n
vf7YvZhmpYejP7qMuzXsmFF5nt3+iClZKN7x3HD0LGfbVwK48B1QXpyCGuI5LN18ambro+4MxyZl
QssD0k77eKMIVfK10Qu5qN53v+MjeEOSwXdDQOIxq9pF46inQyQqlUh+/KccmErpcsDBpM1h5nD+
QkSmjArdb1D04JihIC2wMHOmwJEP+7Axtv9MDEY9uppVaU02fK3lVXB/eO3JTwkC47WL6N9f68ME
XWP/gO+VBseDs/yiysGeQVl0aaNBkBeQuCurpQNOcBgp2mZxiJG/ZjEaEhAwetxanW11xtymyjIh
TSv5KWeAbwctsEnTVvuXOejyehwSg73F1/2u07Mg8tUXAmXipZhxo52E8RdcjNy0XBHzLkb+Oq0i
Qp1DPq5zsLBSiM1g+gIjnICIkgatTEKXN4vfdPim61kGNIfzM/dCs6MU5VxC6BKvLEmt/kchoNWY
C64vjrvW94u634kly8fYn9wCv6xLDOGwWwNXH7b+Vns1pvAQmdiMWzIFimBS4370kTvWmuYEpbXE
wvxm8ADtn0BxIEAPrOVU6v9ULNYQz9J3ReUI+KxhtX/bU+0sul0AX4efQQdowkmwxFsm5yt0Uegh
q6KXGxV5SK/XPSISIAF5hnNLmjhyWZOypXMAAt5BwsJdLGaDNRGMxfbSDBIFoTZOLiVe/aHa1kF6
7aDtFys3E9GF+FwzK+j3CxEGQ1ACM98wSURBtls2ayC2YeWnaFIYIOcZX9QKfi7iH7FXVMEWRY5X
ZJ0l5KVW1VjJZeX+9Os14J3idvDuAe22RNR6vUlwxdlxuXV+SqM9kjJm2CrMGy4iPnyUq22tWSBv
mX5KwidwTCSpcWtEPXG0RZwe2EMjWcH0ptJAsoX9xG2y2hT7YkTev87iOnY5zG1BSAD86fqGOm0I
ZkTGVBcHDN5Uu0FRiiJkIgNU6pqf2/al5fJEg2/0noaSCKvzSU7aVa9clJv6FFnUG00WiMDBREEH
JAi1u+Bqrs45ZdVV/Lz8vVBxWNh43eEonOxYbPgpvC9RrWepNpduy6jUAPdSWwP5NWJ83MFA0pEC
c2aYme3W2rrKgZyWj/vsaVnbf5XS7dv1THkrSA12ANNc4OyVAlEzVhi9+KYrSeVfsYITA1j/wzMm
bWDKObHxy9q2ygH9MUUybXudMnqMTHe9/RjMjFb6dWwotcQIY8BTVvssuANDuTfueQSRjLJn0Jb1
WJenyGykPRWeC80RzppOx35U7qpLKPXeQZ/gviGAKfnJ5rvkSN/VV4L4TbjKQG0ePXtRJtVSStc2
40Fv27ylz4qDXOTNzX5X16Gs8t+XyqYzwfojJJPQNrMM8OF3OlTEvnWMNJands9M/aRMKn6TRgwJ
m7FlBXDCHWOUVcnKDC7Qw8Cesf7Bu2IMffzLLjHUQjPVxYOxGH0WpNk6AeO84A3Rl3nby5jh9D7p
JQWs3OWJ6B5HN004YyEjXDB0jB8XxqcUXnmEqMX3+zgsmPb5Qup+V2syG4sPxIfYVoUy7oJGNsr7
8ekwLHhvpyxIPDkRdiG42xrHnYHJ0lhKqu28MKNjB/KCQb6gnFnsptAxLbnZ56kQtBQxzy5AhifX
Nu7kbKu73oJrDalbTRu/SEad96Oq8TUSQR46dAiYOCLXNZSt3dG4OQXutRcuHIjm/EA8AA94enj3
oG18rV1TwlNYDLmKWOArQrq3rR2FEuOhCJniQVnUxlwpBnHGEJ/p7NIcNa8Rk2sIeYTg9jqp5x05
tJ9FLufMaiDLPx1U5Atq/0eanhB3kxVjFdJlUquGuhiEqyX5jUqAtKEwVMcsD4ct7YxG7njWOgI5
0uJ5n/sLewFLyCXwEKuIClFKyz3BwJJ4PiqF6CI/RSPyAZaBDr11oD55XclS49B/JbranIARuvT1
lTTklfqjIN/MQqYAmy9gHZSGJuBpfYm2NQIhWBhBlhhi9LufKxNB7t9/bZ4H7sVIP1/ljJb5Np8/
yiKIMqMjXaiglM32dU1FHY/ywIQz95G+U32nnGI5Tg4iMW/UnDFyQmMfzzXDGV6/ckNGiOvMD5mB
abZhlHt/lt4HDFFZmBYh6VSeNRrNV3ijOC3LlROmd4nP6RDj5nbKDXd69WK4Hm3UJWVR6jzNsM9p
JjuzTt+JAysUHlWuSMB51U/Kt8cEMEiuVDIyFuveiXX0FeKYEcsTNwIn8nChRGUZYS4dP+1FchTw
UH7QHZHBS5F7xVvYP7mKfAXUs2AhpgsrZ205OH7dmukwEDaME08SYIsHRHJJ20RubYTuRKet1OHt
osFgijmGjM0KKIeSl2McKzN2bowezaWWReMi5Y87TMWgfrZuw4PQhR0o7l/cwzCLTMFRiPxKvbIX
02U7cPUp3GAaT1Q55Xl03k8ee2sQ//bdLNd3qhJXipGijXEk+ZdGeINPzhAL8DL67IdCK6EB68XZ
mX3XSQUDj5Tr9kYnAjR7CNwWb9qQQ9uidqOogEeVwdkxqGhvGk9ih5iQ/9/2VE6eZrNy7UazknuV
c4jAjOzB7PBJq9FRij4SFl9rmJXAs/vXu6KEvDmWolNxA4QDbVeavfPhw0b8YCbZmrRJenG01SF0
nbz1pDvT/6lMpT+cmcc86pJiW7mNI7ZxrGSs8GOMF2J7e1QB7GyActlQlcmG1ms6GKIpkktyQMWA
1ru28xAJJoJg3BlCkJrST5sDEAx6a3M/gR86oaOo6m0UCG6gozNLCCTsMJc3hDokCbd/fjQ26M3w
8xmwF1THDhX9At/vqORz1UMgDRcX4Blpcg98IDt2A1VGVpopMHB7u90pllzFhex/RYSNs2wK4Yb4
lCiATSxjR3ZElEMWlGlTFrQAwzdAWWm6Kt0ZC1g+DtmqbR6nOqdvOJzrdMieEOyuEXLzT4jCogTT
SkvWlqcp00r62CWHjT5zB1I+yBESchE1Lj50GFhBQYqYPnI6ZjdGfGuAjN1isP1zDCigW2hgJWaR
WXWUpZxfhKoKNPH2i/JvT/upKcW0yj1Mff4RexPeHG8LdbNr5eLMGBzL07TQE2DlyP3jPVELWf93
sE6MD8UlGOGoH4Wjqxvm7i7mJEQROJU8CSbsYqdhPdNNikju1zPAuvuwCYITzV3KIDr5P1ph+QTD
5VNSVIJTkQsGiMwCq/bcDN+59Eg+5uJ2o7buE6dqAzRpl33la7oHVAMft5Ip4dymAU8HzR5Ir9eQ
pX8rBChii742tl1nj29ks845i1fyupmZnKgYvBp/Yw2qNO3N/eWCctS5Du6BtBF6HIcBj3J+XkJa
0KawWAoJDcIDIkHkI8eX4eq5z0fVFBTAa3hqj+Nv7UPyRfOJaGgx8PCtyb1R4NthKXiwUrpnBjHs
4TP/lYezt08Af2m2BwsT1iuQHM+o4j67CYKOq315z6rTGUgjxljVyzPwyW4AL7Ww12nC+qU3Weke
RKeSE8R1BTOw5vEMn/zgYEne2eQSbvqvUBN0EtdUCngSorUfnEI8iyW9Ky3mKMojGvmInuqtx0N/
ep60OVk7yRZWn4Wenl/eHLmbEL6GExmy6KyUsPDTWOzkc0uNCMDuZbJvaOywnun/a+8sbLqTZVeq
HyMSAxqPg1doDhZOvpHlmwS4wZDA82IB+8emefmSu9TekejgzVHJm39pcCYYrfME9AUn0jRpO/KC
m6ICQG0KgqxLX4BbsrHfyvNUbKICOThKchmqqCNr4xxfVruyqCvIcXfwsIngrGYreGuuivkXTjTp
rhZJYiStv+FZOxVrVQUWEukBgLJcWF8Cwvl75f5rbhBSP2mzvMnfCGf4qihsyerH6D8Zfy7y3jxW
G63iW1njOHOKh85cA1aGXIR0WKkoBNijUKSs3W0BTKPsUc/QBJpIDXBm0+Voa2R8TgHdIFcqCBxy
v7Qe7FiWy0Ps+J5wOPIFqD7g8snoerNFh6UaqrMQoJ6IDZLQ5CKngjft9WDgrrFLFMMe1D+znq1l
vSP83KYUwR7lP8K4v386fsModMjV7JbFfzCA8szsWwO99yXTySHFoVAgMKJC7EhP5wVOWr6IQU7x
ldxuOunmx+fLB0bHS+vdAs94I6Pjpm4YVx5D81W9tUh3W9js9Ze0yg7cZF345xIu2hPXu32ly+ZQ
1Sz0K2dXeHdo0tQNrxF5INn2ofnojfu4mOzkr36bl/GTF+KsTFBjAYbtGJeqQjGosgQf+1AC9vt0
WZVBTR+E71E3W+apXobrjVHCWVSS8xESIdnhFYyZRynPSiv8vizwqeuFYJRuN525nAseKeEUJzoP
dzE3Vg52WJxV6+8q5RjsNqYaj9eKq0Hs3R+qE6PGOuDXf3vtoCQVSSnRym0Ehrx1KViY17Nq0whS
MOzmByJv1uh6/VDj/sWytoo3VBXjgAz2aeld1YeNYTkbGxf9J6VV5c0ooDVlBFE/6I9hVnpUHway
2aRIQZDDHg5wQWLgWQjqSiRAOc4rv4mQrE3pE4Jzv22S3m83Ujbsr+lGOh9lgesrhqXnewD+fJUn
FkSstFWfZnHbgIQxmKKDGpX/pR0DSitk2JNgoHrxfPwuwoKyhgE5sLabK0yev+Te5I+IRg/pe0a3
9tmXKFqhiNuGDlrEL4rkY78SLInmGTJEx1ITVGEbJSczBHFhHDLzjQgert3teAJDkVbJk+gUBF65
PzWeCHSIFl5mhfelyunZnkSQpwT98j+NEypn7wucvq3RgYV/JAschSeAr9ZT8rNEYf7AbTrEoLVM
lRkZdU47JJ0Yl2gHivSIy1/hZOzEp1sDOl9/cfeyRMLm1eWQDuHSrAxUXNYD1nQzADPekWr0elDR
Cj0YDhO1FgIjV/fkTZ6lSeMYdtAFj4/UzP/AFaMk9eD0QNFibdFdCuB1afU2BqoRFg81kUGOMTma
KISleaY6mTup2+f4gUC8wqRUE0Gb6hBmHHJw8azFZAKCrEQi0k0rO0408twZc6T3Rutsb0d+qiKn
xUGY0UsfnOWSBU8tz4NewzD4tQ6zYpeA1pU8wojW4NQ2Fnrx4lakehSL/+vLWciEmvvtjO0Khno8
lec2EmZh4nSP8CJvOTph3TJexMaYhcYSbWYWuvhfIlOGIgJXsO2flfw3KSx7IaSw7hShXc6vwEYM
HjnyyDEwPFoFN7HJQgICISOUGdjJFHeJ8KM4hIKvwKnF5JhXU6Hk2x+ac5wcpIe3ozUH/0cHtCzo
M06CAgVUq8ucN/+bVy5eQjyZg4cnaQaq05cdEnXzp127vngPvq6a+BJ2wk5Q8oZKxTp2jQOgyE2W
LfE+TlYda1Pif35bY9UaJkqC/B1kzxoTDitEgWl3iAVVVXcvF3OivXNDjSj4XkSGc/CwhutknqbW
DyldM9tREj9vZgEQgDXokx35AawDZpo0fse1+p7CqjvmBmXPyb1CN8anvDMNy9nPEvusznZ0lh0c
Pwzj2pA/tyY8rHGuYAhk18Yb5sf5q8VNbDKs2yo9SD7lryLd1yWnCA5Xv/1X02s+WFI0tDqlmEqH
bKdL/lGMwee3bhCljFhTCsmkSCc6xKZ7nKoS10VM09Ux08irSuqsGsoRymuKvWNsedeA/3GZPui3
jbLuxzaKUexb127lAPAYxGfJmAOVEgCqmqEQbIX9jNTv7fdBUZbxsWylikbKGeBVbzeim/6mNvoX
Z4xanRu3b3blcQsjHs4rWh2l2t0qZA1O8iqIVtKc/+0iLTJt41djTUAvcJNbp7MLRM82Vm3s1TUx
z416GrorNFcvrt1i3ZRXMjx6Kg6NJ+bgXBgBHlGmNJM7L9GCHIi2zLQXzUTT4D0xvs1SpQa/dwLa
rvu/+iAg0TIp3PVCxkSA+mACcjwiOlR7pYynSwufmonsUoTegP3y00eZc4MeuiwPqBIO8WdBS7+A
m4W0l76NGvdBl+koXyt/ivQ8qZXSDTT7IaP6Hiaeb0oy/+84WiLMau4FB08mE3/7pJZlr6DA+wat
94FPFnUHAN3MluRQL5X+sKvcFZhMv4QDkLYP5e9+27zkMxIEXyxL47xkknFNyEEx8kF3gB9Ix4mZ
5prxKnFj9QjgK9U7CwL/QObSWAmaxXE8vVWP9/rdVfXkibRsS7pRB3y4mxbQxIPy+1Z2Tz48veuE
VFxXYg6mjzwgVx1FonFY+oYJMGNiobDxoUwYL/mJ6UcylmklZQE+G8LamNvWCC9A1yNMmPkPXD6a
BK9W2UA6rZpbOZ9OvPnwfDe1cf1FaokZcde4IcTOcSRf2dS4XOmkACCPVcHT7vd1cRFOmW1+8zbv
zP3IIQ89s3v1y0lEAr1ngKPR89UrazN7sCtF6fvVX9SYypVX8ir+5XoKc3gvPa2XuzbUxGIVxh08
UhCNLvGSSa9U5e5rXv4Rq2Fp2AzwB2TgUvMeDI7o670ns7ep9+625AxK3C67R5l7cIbtEX4cuVkM
NvxHQ9qnqDHjAYEkstCf+5wO1FDli1/IGrX2Geo7CDn/QNtf89LqWxSbW9KO2X6SS9QtHZHztr6e
yJ6ZkPKnN6lQE059rxrZQpEBZ4Ci6QYP666qEexRh+aI2IrWjkroi9bTPXRbVBhgj7jOUlziVEOK
cO/jn2m1VFNF46CKtE4BQ5ihCghgVtbb6XZ22lWrSmlcvnWvBJOvu8k5X276lQKycCowO188Mf7w
xKLzg5kA1FrpWQmb1ovLNVeL3av8h27g0ZXA14Xl6sMgyvPdkbWxkpFR9d/fCiQhhL+PQPUaCSL8
WqKmR0N1KXTP6HdAp1Eg8JcCjRvIuk8UmfC0qYls/bB6r994KjzqCF9Nkao5q1ub0vFYAir8qGQq
0aE7upSLThf3SkTJBrDWp5Lbzq4fZ4OndMcwI6Ij/UUCYguvQ/w7ufj27ocJCIP3LE5QlXQHNnWF
TYD4nnHhV/s/z1RYU5I0YLqOirZOa31k71nkJiJN0WHS0n5L73h5bivm6JLAVOsyyx2DWyBy0jsq
p0BZB/2UBYm/D2lgDzWrtRJwb9cHryhQOGUzv64XUsvw+ro37qDzweP2IBV7KXCrW1RVEGP2ghWW
oXVkKEWq5yIsaQAp1XzwtKB7Sl7uRFHQm7zwuuvfTkVh3Z477t77sEQPhGDnWmzmuzsPpB5AVy0d
8904ml2rJIT5p27jwv+ZL5d29igU8VrdDUSmFvBztj6GRRYFMeno8o+oUfO+0UT2E27nYQHSBMQX
fPXjMl16GQvPYyfonmc12aGNAtpKbKEsRfJCzB0Fn50WBDe2Vliy/fg1KDAIdVy2pLp5AkOf1UAt
iXzR8/Fy6KdJngCUTI8JpY/iUqO56GkIL2L1BX7v8gmbzQqYhoB00L8O8jDCozapi1ecUJVZkGEZ
mq8xeMU6IFAdUQByiO79opTjRo3Rvi5V/PvQxWtQO1XrNRVsrSKNVcOHRezTv6wzwQ/Rc+mtAocn
lMM86n75PbWSNapcd3Kdh7UzubeM8yB71mlcfgMCJ8bLKW1wnOksmOjPSwgSGssqp7JA0AOgoe5n
SOQuZFl/grNgkMAQlIDC2e/OD622xO5xyZLsyF3uEMEN9MXu1QUIB0P9PxhIAurR3U/xNK1EKjS9
SicR5VT6OTR/93a74XYuS9KnL4AdyZg4D7TVCqwCMZQgKN30scGmxiZJXU8PjMN8CiS3oFRnHHi7
IJDtbli8NTVztRruKWfTqSKMe900KPYcuIEuIRO1RXUdw09iVW9cVLsZuEPeRX8YZIHdgu+LGZ6X
Kp9Zgz0YCPDwZWb+AN/3VZ/zuPOWW8Z/wCvT7CfT2ummmcPONKP8AG0eeIXRk4ec6tnhwe1/dW9u
izfLjVce358ft7wR7idreoZJLSD9uneV6JxwQ9WrGxsRzE8IwKsUCClFjpoqRazy0FXMgESMt9cY
po9/xQWbPYjN8gFYo7lB+52rdyQe/w2BjHQqqJg0AaQtdIbJwiqlg+W+tlebALbPE50DxE1pAmDg
PVAzWgTTSSrJKgDoI0Mjjytn32DMeuhXWmY/2KjoZ0X1Vw925PhLUDt+QjvycFjM1ChPIEiejvGn
w7XLFa9aIsxKM0nnQvJbLlpSs27rpBJ6F98eXBDCiepGrCFA0r6PcgODVcAMl/7G0KX4wiNhI63q
zFOoeq8woW9y4aOn9Q9GCEbOUCq60pn7Z5CHKqLjsgwybjndx7M+GUpt2tRLmlGWGkAUt5tLlxMY
QPkGkySrCBNCLl6NStJr7QpbAfWSkUkgRM1yxy4hC9KqXOXezRAxnpS8okwrSNHxHUR8D+lE4RNb
A+5IeLe0mBfMe3hqOdbACrspEZ++7kM943bI++1tfRleLqhQ5WC5ZZmOkuLt4eqyG2Cam6eeqW2x
YmtsiCRucedrPTDtANBPQHYYjzn2NQScV/otaTdH4CM1qcp2YFdArDQty15OXfdG9i9mdXWBKk1E
LNbOC7XbNhyqh+rkxX5G7+kl25ItD2iQXHxwHVpmGiorUZF0e7MAhs8cdsuZMZ+fCzAKCFeJqkEO
6iUh0OSJzk41xpY0YWkBOkd7YRLqjqb5apHKZKCa2FHr9o97r/oHiJg3Xzd61Thps3l13ys6+ka0
7U6IHa/MPNiq2QtpvNvCIMFzzAdyXaxj6DKLMM5ulFBab2/sfuBP7GeuDkmw+uQyA7qQNWVI69JA
I4c11/kdSC4xwziA4pLuvTRl9fFoTt6Sdq7n4zgUikJ6tfWkTY42XlL4jiLsrA3LQz+Vbi+bksvV
3ZHIVtraK+l5bAUQJyx9144Sky+RBR2AtT7rrpLJR6Rq8wmqONhwGAFp3wW2aRWs77ukuUraZpze
i94SW45wBOeu5xygzsLk3BMmTtrECe11Mv/cBHokBQ4+UbuMAphQRGetpU35Bcx9EduMdtFFeFgP
9b7TQ0ILsxFR0+vM/hXysmt3fy8ox+VNxrH9mAe2EvxSKb+jg+6VTnD5Y6uYOG2BGZYaqaD3eV2g
FzVO8CJs7xiLW4Ul6el4Hs956rX7ebZik6+gxQ/4FJ1wmoVAYw/ycRhShBtZTaZBnNKHsvIK/CHz
0Pn5tPfCbhwS1/bWciCHTo9P/t0Hjjbw5qWkEVIRtFUnoq2yzxpABGovVFR8GL5C14pyem64mKO7
stI6z0zvFqfU9fp/tY3BfzrLRRTTU+lxnvi3clX/vdW9y1pSGj499aVAirgaHLb2UWsKU/WZ3mxJ
13X8bH5dI5MDnxgKaxqaBNNkSKL3EK9ZAtpPUjyAAb1UR8D4yRuxG0YZNLjG973XEmzLd/T/fQVS
9LFv48tDgvaZd/YqCIkdMMvWY1L3CwdjWdC7FUio6ow/s9R+lQ8YclESHi5z6A82XNGJKXbLyfRo
Ryh5PtEsFkEyQKF6dlVo9PqqmjRsx7mSlYtq6XPzfic9obWkvjOZ6vRzzZSPxHOj04tomV6YrPaM
siT3/5Gkq1fjaJBjdFdI+ppjLrrCMIfCgh40wVn5XVw8i2kmaFWYud6DE+m3w+zYsDxeiGZGmWod
nkv+fUNwfSQleKP2mvMEKiHpLK1XR//x8gs8fMQbcr+fG7UiI74+nquUCbDsSYU+XcOowzY3PJDE
xUx2wshSjg7FcviBBicM1jp7kaDkQiI8ouEQ70vy1cremHKsUDif4ou7q5H1xa4We891KNBWJNGd
bPldLNv9kpIoxX4A65nKnYRzfk6YBB45IHgU8R1uj+F1MI6Z3h++n/U7U3fTWTq4qbFTba2Ke8qE
r1WESjpvu2FGTB4LQDUIolMD8IsNYWlCVluhbWS/Pu2Q83X+G/f6zNUwALBSWOsr9Nb8I1LVyFj0
XFLQ++wlS7JWiK1HmfrGj9DklExlLUcpwmVe770AqIcgWWJm53dZFsMn+dZPOgUswN/ldvG4NMbA
FETWkwA4fgMfoUWyaebco25huDGC/HvLreRbNnXyb3aMh8RYEcr689/T21yVV6XFuYwxDd08KvKj
4hHZJvgg73ljmwWsjQvwjI+AQsTINcCpIQAyicfdDTvjcC0NqMHwSQ2f9kznnmTc5h7iyv/GTRO1
ieRUg9BBTnTeEC3nV3iccRBgV24U6yPc+WzE0aBAu+nFEFB12pDWZYyscTLQKZ7QbxL0jIGylLaL
+1ks5hyQIz069AjSHEMonStkGAvnBaDgvdo+MzkqaGBgVepTsoShEAcqf9UJ9zKe3eUHkrxpB5pq
1u0mzli4s0WkMCKcOJhhfFflonEzjoZdZLiIAu6K8Vb8VcY6MO5gUqQi+JOPL1llaoH/LT24J4w1
Nwlzzz9MMMbfrr/yHHXh5n9QfeC40yeGif6/x07/zSxmxNSK3UMAosXu1rB08vRvxejgi/F9Iwu7
qJvkoUeNvKQ1Gs7T8kLsQg8b5rvEjIRolWdXtiqm5E3bjkZk+heayQKH7S2FI2oF4PlRLKgsjHbh
KWNmPpB7G0gjZlm84Du39ugyPuqjS3gUxfBQhS5WUvnrjQ+PsywbuExBs+gSiWBMZ2a5jwSw9C0H
X03eZzH0k3uxFgdDluK8kZGplQcCyLOTaAyTXSZ6TYembCPCresKyIhMiN14optH/Y757y5QKopI
hFk9aZNGeyxunAd0+G3YkWOJuhh8Qr/dtDI4jxXPhkJUA901NXbx6K9jOdqhgIxJ9s0y+G/t/BnD
Xx6SmInETbuG3ohnT2dZ5lrqMSPkmujkZGoaqMjbG2ZMne8fP3TIdbdfxfgOFZTY69tT+YIDJnAK
Cpp3JjsQxnbmu/zbm6kEhW8oODdYNuBKBPjLUBmdxl8Iesl5w9+TKAkg9qMIHEf15NMQ6vNKxc+X
DzZRIOxtNjhI5POVROUyn5jHGUxkOElt19mLFMYTmKn3+AGd5yNw7praUBzIt0uBYR1e7kfPQ4ug
C+NPibJ6D4hmT9hQEZQHKDQpQtURxw3De6A+A8D7tLrvTo2D2ILZX9ZQ7acT/JiVTDCsmJ6SYxCK
4oBNlUzHDpqGHwWNQxhAdZatqppuySa885MFzpWw7KQFB2VLL+ZjtDAwgW1y/CHqCEob/QdcIAwZ
gNmvSgME06HVHouPGG7u1Ldk+3l+NOs/DY85348uKnRNh1nBdI5uvA9K7K5IGXYvCOgaBWO9bhMd
RNfnlva0AOneE7KRh00TYCX4+lWx9a2EliSYo3y/u+s/mjBprFSCggRf4Fnqsfo3ME1CoLczLYyL
iWBjNPg+2dwf2MLsrsAd/Vt4Tn9ZSl9l7E/a4L+HYQERCUCWW5vR/qfl7K3W33kzmujQTAIoAp9t
zjO/zikzc+lfJg+xqRRiiXcW315EleC3/uSNWCrkyALRHqgoWcOIC5k0CR8d+RHOBcvHZqQKOYOK
oPrsuUOkdHTnXQyNAxbJGiGWh0FvuGIa4gQTDn5XnBkmhTit2FwfEP3fmuvyo1P9NAKKxyv8cGFV
Q1I20kO/RgmDU5VVys8F42+o8QaLGoBen+SbwmVnB3/mDz2jSUylSQ1Yeig0b4H8FCdkJ8Qnpb9V
XB0lC8fCIdGzkbmKqTIZgfO/wpKZDno0reSw5HPBiNgyke4A1kDoTg4cCYPS4ju6Ms3DMCjinLb9
tqfJ78Zir6u2ak1BMGpm7+kOIeqIYCcwUX3+Q6JIlWrh4mCp67iIzyhBz8lUzlGQRGwZ9C6XCf9q
Dcw9rUYILHdgJPiUL3OiVZHTg2glo6VX58PyXYq9GqGdpn8Gu9WDv/xTMfcbi8xFvVDxfwltmoYf
qweBXEIjKl9HMXUw9P3y8TVaCFl+sV/1DTSboxImE5WspHDMgxdRkESt+GECOJzJAzKf/SXxMrFK
XKlDu7eZPiW2JQjnrmODuMWd3vJ9ERkmOnjKCRdpCWTq8CrTfwekKlVTmkF6EbbuVgwUClemVj84
mNetYKKotbdDU5tIDVe9KVu/p0ZeDFMSAxtXqZtNMkFrojxQ9Ba17VkjIXJPLuo6d/0Sy6KYCMtx
iMG5ckWKfgTo0m9Ddlt8LcpIc5tFaPjaLnpQx0zmR2+3/5NxSqscbfMPsXqh7BWLlciOqs3MQS1/
3hI0+e1RxPtZG4ISRoYyErHJeFL3JXxr5B6bh6/Y9CqpuHrwT7heYfGH/00PHADNneESP9TAsR+U
9d4vmzNULO2swCv+2MmNaWZuB6gs2HxuQRf8DfKsgVCwop3qYZ7wvC5kVTnEbkkPF5wpIESugHdN
OlpTH2p5OCZT8Rm0NKzxtaNuRR908Sm9uDAv46hdCDgjJS/W2T/e305Rnu9m4SF66YQHRcZcHiD3
sKiUjEY64d2okpY22OCVDetDLqHAdVkHL5VVM8Eu2gPrq4DuNvt8LtlmwIJUaKU9HNorTOaLNBjk
hf8cjmBnVk00aGfq11C2QYq3p/QPJSVUlHu9i1bt4smxoARYma9o3ndOypomTin3mVCYcxX8OnuE
/aXd5tiqx8UdH11AJEHOJeYScB1lvb9rvByYIR/hPCRa056LZzJgLuRow1WP5vOyslPIm7t63aol
ykU5NKA2UrisRxJl4LQ6OMyJXC0OcXzdlqSMuMcYZCLW++ReIhVE4YeC6wS7YhiAh3R8yanuaXYP
9CaIBBIKyLkKdZnecxicYBthID1I94UJeT5xZT0RCtVPzx4ghc9ncv8V0FhuhebPcX9stIJ48/Q0
nXcO93zxMeFZ9KY0wkDxug5DMPLb6bphQp8sdUe8NF3EDzqR6UEnnJkulIVq5Gr5SWn5UxKvJWcu
09rl9ulobZoIwB85u/Lbk1Cjws3fQTcbPH9VwZzv9o96IBLT6pCsxjyzWeO9sQRcnHqSJDHrkCDB
XuMkBTrfE7x+Fo1+rNTfKYaaXUOb7DT2uk4qYtWqHs9an6W0ic4gGWek8ZhYv7AT/jZBmC6MnviQ
Vol7SfZNB9r3LtdFlYirdXQIlPrq+y8yGUT/Ypi2JYUVwYy1Q+ODpf4YOyxlXra7lqUKfTSJ3YSL
qXp6cs6uqO7x2g0nrTO8vRvKlN36RQE+2yFtr1FbQKsUloguIdgXWHPfi4gH/1OjYmFBTVr5U3zn
uq+2d/aBqCGX9oT9247n+YXGDsJZvZvwwiOXa/kslqg+MNZKecZgJe7QoEvQZgSlcLX6d/q8kgY6
k9eHRiVX96dsoKw3BWnslbSXe+EYT62MYzZ166LQGw5o61ch/1oOuw/zttvt7o1RiShkcFr9oQAZ
SkCKvBY1vL3S/5v/qcDXCN8FJdNAAMqv4KL9rEdDon0C9bkZiNSN6o44IHUEvzLciKwt8YX7QZzT
UdhiAo24yMWPhmMt/fyxd6JqOuBppCvn/l1D8vUzy2s6F9WeXmLWkmNxWra131hsbvwXKZEwMq/e
NXXeoOgp5xglDAdhS1T5bO9C+xz85/FYldCftxWjAF7tuXOxRWhMwWrzEg62k8WI2LWLHJdOp8BY
NI11/FmI45ukEeC+Wo3sMaso0aVct8gVQAkmwoRgD82T7PD+cVFjVf9fK7QancpI29mUQG9ZDkD9
MUez4Hn0cUDgmJI5LrQHMsQEMto3NqWGQEF9CTtieqPbZ+keP6DNwKbn5nfREOgJPtWHNgKLMWjZ
Gb5l8aN9fZb4IEta8aGya7Lh8CI21TseePfxKGklpA/b584pM+M8rWEDndzhR6vs5tHNa+dCC8tw
PxpLQXtRff7GHgDH6EaqMHboNv3uHxxnwCVJvFsikD4+tDx20wgJGwgdEuzZel9pJVAWzNvqdVmN
FeDTPHDkBVJlkanNzmrSbXSVIlxusZmxP9QxsX7UiXIKANaoYvaeDyL/ZVpFcjlYRnnX3mRSj18p
6b5+eG32npX16c0wGS6BPaGfmGi7vROSuF6mMEqakG7X0g0pNXNiIw2WUY9RJCEMi74tTFhqxEjK
j6Fi7pN+gK4LeHlWV3Xl/Oh8ddSAHhIC5Uos2ygByF5fQzvbVYciKDz/4otdX2V3ruaPwFOyZ0XZ
GtMB9KgjM7E3iJnVa/c6gG7b+UaOuO93Nr4YuJvvaHRX6VeJ/Ty1dMuIc0b73aTHDW9y06e29zZa
mxoFwGZ8AlDjWczBlhGOVQ0AgXU8i4vYHR/6D80FSRbKF7mLutj0K5EKxd9WFF7JiL2tWIY5sY4o
+WYsvSt45KYMScCcLTQYl9u3moOxDjRUgXm7zbxOjNlBJVEpQEH6BahPoVFTDC/aCLJhcs/ib9l4
qDbiV6zDQIuR81QdYd+6ndsVUqCZu3vTWe0eVSXCpI75WLtatzcuUoDZ6kC204gM0AieDqptqZ4h
0rlhaPYdJVyAVItYezTjrOoYejb8lBIIrAc5oG3LMgRJh0hppzQrr1EHEPRQUZ07b9d0Osgt5Kw7
sVBRfL4g7ujmjmxCYUNQ7/YVR7PhEXoypadwg9eo6UwiwYP0HWEhwu4TDwKyNga2R8aSiFcG/byD
vLQ7vyyj1N5JNLnRg72/wAxRX2+gs/OL3R0b8GbJBkj671Y6r5AjkSPRg8yWa4V+agD5Ii7dC7ch
SUK4LESld00V4K07V0W6Mmqhx3s5AClMtdL89Ou/+dc4WbNGh4GTVFvG+9zALFcj4dyxKGZG4kcq
SIm0A7Y/+6e9WL94nMoRMCblih0XaGKxTQ9616RSaGSSMhPd1JSBV2VYBIq/fVd0dRk76uN+7b67
Xa/swSRPjob/1WNd8fUMvlySGZWWoYDiL32BgyDJFLCRwnJtSjfJqAT388+GpbSqXLulkegXt8ah
Qdqt5F5YJtGgojz9aK5w1a2QiemJs5TwS15EykoRHt1MuroBb7mzl5h8iwOoyMyY3Yf2NIQmXAkE
0v928FM/icCNRIiJoJjWyDDnFszDOC6GSBQNABYnBLBM1MPgTxGcMKHs7XlfzdS01GFlaIbCCFmQ
YGYefhI49VKbM5fcfoZevfJ40LZ8cuttZAXxYCM/SlbX+/zgLtwK69mecvpbhhc3xiLCmANw4d9i
82xgA3ShxzQp3FbPhSStzZxcL4CT0+M/r2/uqtq7KROQCGTvb1xrk8zwkv6zJlHbxKlFsG+7uU2z
HQJBzLXJ3b5DgkRAJGbVJU8Jvz5tNFVBXZ6z5wWFOOTHKcyhw79UMQVWhhQiUDdrCOiabC+uSmxG
BWeAjLvfncj5EV5PpFhJ0glJJ3a7t0cvDURvwipjaQNw2cD+F5Av75aXNIelzP1TKQXSUh0oDkY0
24u4utfOOIb6JEli/O/s09QFTkhRAg7Z+P2/q/o/zlKg2bkwozy7RhIVlxrMLvJf3w0mmKP2ZIUP
vb+tNgXzvpWyyotm/0hmvVglt7sEBpY+QBkzlZ1hD+U0K3y3hDwJ6nlnk0B2/S27hfE6MesLe6lZ
v6TmAMN9IT2fA4MsFuKQKtX+sb137Wx8RYtFqc777We1bnvMxOD2KUOlUXsQPZlYk1Wn3OUWcif8
fkNB+amm/U9qb8BIgldLztA4sNbAV7qkug5lAmpjnVyQ6Rt3LkmhIJnPt44R+kse+ixIEBO5xsFA
hXZQpPHuLiAyhFxXhAYY16vi1rCDK1yynrH7DKC0m/1sRY74OFGLKEDP1I0gfp41rAMcytgqEoha
n0+MaJ0cfn0rks1uhy6i7Hh7zuwkf/sXgujVcPsns3Hq0Ag0VzAWnkppGAiScDw18OSPC4lhAFGr
CmWLtDOpWM4fs2cEQmyA6vhAUdfaCLSiCaYp4E0aCUfIz++l3XJzSgy5uJlxj+PczcVnomiTZYgK
zyESkROTdmvImEoEYKdDsuQpnh9A9s5d6hDxqRuC/5LoaW3+ikDx9jn1g6/SzpW3P9z19HECrwXc
C/IZRPCq8I1Zc9MR5WX0MYp6hcH1TVjHOOIVNJil+KphiEr+95Wi2HCMzMYQyZI76ooacumiP/+m
/ZT2Tbd3Ijzio0jX/0KBINzr11XOYqAXJJlzmr6sBkQEocDShPacla8NQNZlVak/RMS8d3xDlW7U
mCD/hIJ+T05JwOMxi/h38NQfPknRjulkH5IkE038XtLS5hSukRNGr6EWhI0tYYDCrI347MSuQJh/
cXMqfN8JB9lNT5pCQzB5d8x6aSoTMXVmFYxsu8BIDEJQ/9REgTSO71VZcVHz48yOamTY1nyr8NW9
dMVidQkt4bibBTctdRVqY2fSlTOWtiA8bCi6L/oZZKmommGTJYNvOMtnzpk88Sgt+/S7+gNkI+c1
XI7c3TdqluoNnd27cdp54TW0qScwMjL2Sw16zFmgvVKab96mifTq3yhX5QURK1Us4XKPSgOr87xy
tc7qYIdf+Y6mWade0QSQfuc1jTTZ+77hbFg1deSG8/asu3O5O7lLipAdKL7ipRsCN5oMCNo+JIHd
RAFiqNwEkU9BtupK5oQ58WexRiaCuQniBFKVh3wAnAoIuNhJW7uRvLCf8/HHUXPpBUayUTmHVDN5
A0lvTjByu5NyOw7k3IW61fOe8YkpQHSJJAgslKXmX+SFXi4hunq9Md47j729Y749ViN95bsFvkKM
wv5uq12eWAEktU1krBDmUTSdnymK6N/O965Qg3987Pwg921y5AOvhKj2WmX378/L4ZeYiluMh3kx
rn5Lqi9p1a6PcvQnqmfwJ++sxBifpbvloyWriH27b8/JVk67Wj0gzcMCrVyoPEiqtsWSNBSTA5Sd
jR9Mwsv6Zw4k2197UD+04W7PWxNQtX/fQT2Pj1FNa3fX3iUI6X63RQDcocC3aYz5Ai3YRlnqnsND
q+Z44pZkLcqr0Z8kJ+cgwqdFoEqWBA14svKCWWMF/9C9sKNLO8KQw7dU8E071vrM53/j4QlDACxF
hx4pXy3T5eoP0RhQ6QBzylGSHaV5KdfGYscRttDCDDXyx3rW7Opwb4ty7wXeZcEqE5dDizZjFN9B
/7VUdvbAC7vqO1L8bJc/luOU332EHQm273Mc97NMhcILEiXo8TKEP5TqHxpmauiCBaddtlhqguHv
DqG75M+j1FgKgjQEbQKusczW+lEDK5jhJxvcan6LEtHuNW9RSD8UmAVXsSl8us1LuAKbYeNWiTEA
Ev+HNejt9jIT6wxMw09aaumxKKywxqkPdGGGlxGZeLiyrYQZHooS5imxFVAdLzMVXEP2/FAbPmdG
OMJy98oOXilb4JV3BN60eOSneubwWsSs2ZaKeXrumn+jtlwpiV9SEoaN8XIFI12lrw7XcT7CurvN
i9vp64KdAhsMq1LgR2xz35aHc1ERqBW7vVyUmDlP+3XY2C12QFAL6tp3t9Y9zIKiU7C0xfLwQTRQ
BwbLDy59K2FGoRPMjnCNMbyeTudI8nQHPbl86LOtgR/YrNVD01hm8ktN2VX33YcK2HFQngnRhkNG
EeWuiAVNWBayyOLJIjgnE+sAVpbfDZpnwNLAVv6exZoVJqJQBtdkpf47etBTo1ZpKOwwXu6zB26s
Rc8ZG6C6jIB66GCjMi5GPEhDK0jD8j58f9l5MfMFCwfEEQCpg8J/0e9JSNBFdNNOPzc+vjK6JWeL
Ss9boyRko3ly5XSA0RlAYNPqBdoqVNgH3qKRubbQwKBiWwTQZp3P/9hgkq7TtRKBbkJBbcHpOV6/
X/zs1rR+q26h/aus7CK8PxH4IvNQ7obQZCtdIFPY11P080yDtSX4i+z3zOMPFFYJ8iwygw+P+QSI
fUZ1I7msoPPNJg712JjhjWIoMXFsJlZ4ga93cc9jKS1B4zMDm9eYaz/rQL+9oY3Ojhn2LUPsHRXL
DPxAoQxYS1/f6KWhaut7OjznXsHD6oJatiVBR6GfJuJDj+HcrKV2wAuEuka7SiojCb2T+9XgJYYI
3mVOU6mBc39/Oca8sDMYMJ0wAOkEBw4+b5Hm/5smvshobeyzsKq2Ovl2eBAFT/LdQDFdlZQ3EbRA
E42E337Ew0NV0Jd0DRQzI1zPh4vrqUt77mr4OcLUhS09XKU9bUHyzaV0EqORrpzJTPV2bQUTGbTJ
dpkxFjGnw3lcthKP8JU4VCwIszIwA2R9PXK92o6T/D+wOxQQBa8g9YXA/P1qBlwGML+BkBDBkirm
F3viQ324qgyNAPA0XOliv1R5ubQMiYf+us5RCgSzv+IngiuBPg/yHBUIbqFx7gvTCQneWBVub6vU
hmKcqyN6ypGyDAIqiDbww/sfgXrGMGh15xJSvfBksj6bMQij13TCdZWGZDEyUr039qcik67mHUnT
f4fQeYTbtGVOIkY9GMzNU3hHbwg8xSIwp/PlpIJl86RcO9VoFN0sxJ8lPv4VtwCtbk/gsceCpdA4
6OMK7UAeTdXlXo9HGzNQ6fO+pK2w06zPRP4VFyee+F6uKSQHEL6YWQwH7uVtOdedVBpCqpfOW7Y5
MW7brt0C9B5+Xi6XAhPdEOzpSZ8Vs9AvfHhbxRftcFdaFnBqVVI3bbkM1rVBvbLte757WzbvXIvW
Dc1Hd2VPi2R7RnyPjlrgfThcGiCDNjkjELDd/PrUVuVR2Pk3JAozu0NqQGl3nWM9tYgyGfyxfgv5
dw4j0dXoHEy49Mid3so9fcFdke2sHl1vdbawD4oB/aEbyCI1ER3sdynfmmvq16/1cAi+BaQVS0CV
vF1ANAMGD/HcU2j6KzURw/u1gWkheKNG3FPHCaoXSqvxUEKKLaLHRFiEAai352VJVs30TSTCjYSZ
JLDwTvBnC2854ky/mK329da0EYVOZIoWWCGG33JtUDUZLiABZDOuzAJtUwVvEv8lusbjO09wAWWw
QugpEbWBaWLm2vcpA87zs181Fp/3je9zQPWxUQMCMRcRpckXi/3fdoL+HpZSTXO37buZ2PhTq6XR
QQvvOzp0QrZvRZseM/nVzgpOG1cCt0hof2MfFE3M3RKdtJiVLYbJtBE36S0ClPQ7l99iAKQTnWjP
+v90aqCYvUH9aQsLT54JBVqLckGknLWAm05ztb+MXQKS2gKp1EjqAqVVvjbm0LB8KF0R6SRWkRvY
xgJr9aB1FXvIUYLLvzXQZM3saadOnPe3YzVCjob+GxIU7nqKtFNYZ1gEEX4PUgLpE7C41vWuGb77
dU6fNBC1tZQ+MDC+f38L2ASyzKow0MucFwNmcifwVRqxqtZ7T5qxUj6Q0/5dQ6khgHrhzKNHovx/
0wR43fS4o5E69dkgADbqrwdWzTJRpwzLMsGrXmZHyDM8MfBgeXVD31GP0mA9FU0nlRXsqZpO57pi
vdswJFEiRgOGMcc8SO8XCSAZPw+iPUFRYk5qtwesqowKOQ/8bdLP6qFthoNdY3Msu2GpPoRNSDol
YOJmx6rNuDJ2ModEYcbbe26lRmcOWtjGiGfFpVb3GpPU/oWnTEK5vpyJB8VfOfHQP7u3ivu7mnnC
Qo1np4VVzD4vVq3fStUX1tJlSHY4b1jClAfpgBst5jMxZRlJRD7BIV9nlXnL/4FIkw82t9OvlDbz
TaefZRxHUodhxeItOz7gFji/k3CwHuqPWd76CQ2Nc6Vn8P65dnu+fpRNzvQdjnAebw0BOP5FA3Dg
5+ClZu3TMCxHHeVTuNk4QatdUh4vANF8qn5FZSuttJHYtTZuRfhlfxAQxXWolbJZl9VNOLpqABde
M8WWlMrgxTgnF76isSD0+8nhbAj3myvKersdHn0CHYVbMhy4pglaurmNbyak6xpf7YtnKzT4BAUT
1pd0OYNCk3HFmzwLNWzSPvOORjg0SwU2eceJnP7OHaiNsdk1Pc9pCH0A+C7WR94AIHjl8FAb3sY+
JSPj+5eshaP+NtSDOYJrDcWs1wGSXWGy3/9QQ2jiYTr8ziULo3pIEkMS4Cy728keFSZWULbaS9+4
dOmTOX8kSyTqLMQ9b06XvGLU6JEgYYSMxtlZGOS4XjIu8sUS53ypmnMSWVpnV/ZEHmH04PEnD6r5
zWRGSzy2im6caFY7GxGRwR61I5g/h1aDVZBnOk7wk8WCgzjVoGJFlQfvsZ2iq2D5ramTrLOPWt4/
xH3O6yaTSjlmld/wQdlrHXTqkkZ+OuOKVrTZHngg20uoWSlb2EA/akPlvwZDSvTElVSZta4n422a
9HSNXkKnm096r+ZpqdhfLZBD7Ax7H/ZvOEoQZVHBwG8vYAro1bTUutngZ5quE+t2MGYc4QiMQRK/
qCYaj+/LW1zu3obs07udjk5IxdFOnew/9aKjXBOJw/+PxnuEdYOW/x009AzEnG6eCmnhVyhbWsOT
A1wqb2CH6DZ2o/s/sDs23WuoXJz+TgpbkShnisirzWLqHRgcx6149nMY6OmxJVAE50V8y0AX2MFG
jwTh5mQMlJZwCYFZQcdFqVsscykC07sROjTjv0nK9cyA43/fzM5nwAs2feFW6t/9J8gK4w4BZu8C
KsoAGoTEFoqUYIIfDZzWEGrsXuHhAwz0aBn+UdYRW0/TcGNMyBptJHYz5XXHPG1vvkri6nIYfCN2
0J7kPIM4Iia1nBqKGOjUvtocgEgIuZhnyCsIDTRzyh33b5SdsRSuHFb+GQ3EZxTN5AhCIqa04pI+
qWRYDzJfd56gLhS3eJvLvdWiqaj7UkLFM8VgjYpDGiwinmMmTZxev28mLenXk5NH/i9MuH9vYA/7
rXPXsEbQOjQu4R/YSpD/9t+k4gMD2m2ghN/TGWOICPKdeZET4lQojpV/b1qS7ddyprjIlHt33Eap
KGeeIQFVqfSeEAGV+oBLshxQY+uSgwKfjakeQWsi2sy6bq8dHtY3pvtk2dFNacwxnWQt9Xrfgoft
kRGl41ZVwvQIK7HgIQazUk/0nsDVtaaiw43KPjJgzT7TPPDCeKmXJ/URdSVXHquH/oC0elj8B3no
JkrdkKV35NRS9sXvSA8dm3hixFy/ZMYzJKwsB92NhE2fLOi4SxBfLN23CnA2q3MC0PDof5IBG57K
L1HXzVilCOOQeztywxJoRFKGr3tjgjkwx4VEDjZ+UvNI78te4PUV/dJfQaL9wgqfUVZX8FBLz/+1
+2TpZDJN0nmKUzobdk6we4dWSla075LTxjBRdBtQGF9uDkjou31+gNuhoFmbZ0eNLp5INH1H9HV+
hTeF8GVjHGutj2gbjW86y/phlyiOL7Bx3ZsmliTiw6CHxwnMyh0R9kuv+sBMKSoxz2MMI5JSpvx4
2R2SsgXB7c/WK/0/f0lYIEdUbPU3OqlS2cBcHoH7owlcUCtTJoIkVhpkoRZMzyJjWHpCjQJVks8c
3dxh5togjEBQaYHE34Xd2h4X6jTDqHVgHuVrRXNFe49PXkK/uuq6I2C2O6ACA4XbEiOsJKvvdvAY
u9X8/HfCZhuWV6nygdWMW0V4Sdg5vKAMAh0YdTrFUmz1ZJ90/NzM8uu0mSzfws4UGDwf/dapEtd5
gJSTC/tvnXRtNUF+QloGZjzEftvdoJch/PDBADxiqiH8s9pNwefXc/Dmf4Ai3aLC+iC8vhDP9Q1G
xlJJNw3AePE/1n5enjJDMizEWxj2BKoo5K5d8CUEC2SoXi6rXbEMAKOwOueP45A2nZvLnBoK5Wcg
MCxEvFFdpLYdWQZbaLG3xTqElxpVj+D9IJoa8aL7Z+FY0RBWS1Av8ejArTGX5EnVO1OnECSLySXL
1DA6CKd0xgSoUwzrh+sAapPeaMHY9MosCKS0uqW29QRURYhmuZ7IuaFW6CnoJQ47Q0cpzXHJcYyJ
IIV9MjebwvPtFBkTYYfaNSr2cCO5Uh4pqKnz3CpU1vU7uAbeLM8R2W2peRBm5t4+O67npRAJeM3k
XbZNsZsalv9ciAQDy7GYp75kC3lQa8TB+9lbr10i/ODAt8uJKvdPjEgB88b11toxRAkrPf4mH7+l
3+fFWoJ8rskXcNxGwdSyGdTeJnQcCgb2Ttw5K0ne0A7xiN+eTqSDnEdbGvlAPGTyIZUBlMBhGwBW
GriaRn1K/1z8PBtOOM0t6HpX2n5v8+K8nlKxhp48/9kYbvRnxes3e1191nrukeHlyTBoicuWk39y
0FdOvOVe6OigV5gB3p4SvvR1NavGMBHevEB9phdf2k4iRdS+TSqwwLP6LE0nXJ/S/IcGlHLNXFNQ
ncW2ZpdJPd/jXuTsuN68NumUsZpWW8vs3c7pPgjsxyYzVpoczMQphPivTjfBN7dY3LxuXCXbjrfg
wEtaoNUuYPilLxxQOc4UNvLlfCGDX3udWJRlpSa/cfcHthe6oYdH6a+uwHwkgbsxJAdrYm0Aq8u+
HpFjvYntlGMpmhjgW/yEowqV1AU5KkZCtzp3+0QD6bMHzbWEY0XDIAPPbv5BKNgb34HIEvioAjV4
EwSlH4RTqhe1va0G2DTsAQmQWt12MrneGG7HV9dMgHgLVhfCjGY/rOnF2gj6cZ2Cp6bjopXwamtn
H2bjpniU4b4Vi4ezeggBK9KDe9AYI7cZnd0mqJyXxFjWG9rrVoG4mj6LPlxpWOG1HxCYksYcGi0t
TB/GFpVDcbMrykhjPcwg0+dedvHz2PgXPhq+6umVUV1nxyYYNjMJbdFzTeikvXRyZIzze5PJUUAS
lAmApxqrqJu2Sg1lGLrOpXQ4oqcB1xu2J8VR0aaRJJBnuPUH33KhdF2dJJo//Eu2NPh55J3+zG4F
Xs5MbUc78gtlarz6Bq9I3Ul+FMnJiWAhBdHRdq+CttOJ/1F0oHFxw73ydrtSZismZm/YYmF7fVea
Rh98MKkKvOLoauWdLmzZl3/lbmi1e79xmiIqXDaMT0ESskIZbACyIZujqxB2R4rEsJ0HwaYKtGI8
lYnHeb3oX9S+2n1xCzLo9Vm4w7BI0u6nWndcNePdWMrtNOumSIwKKrJwfHigrQaTGZAqHTPKdNgz
QFA0vr7/VBGeELuuutU1c4YkSer/taUbJA952pNit3fDqdqOcYdFTX5nAbjJSyKVJwdwWy/DD3On
YtCnJBrapgEdZwzvcsO98+EpA06licVLDhuAuifkMyh3NFZChqkHOnicUw2Zy6GHd8I5ZRwZy3MX
HyFvyuDtBfgYFzR4jKKpWUJxcWfOg5A88eOOi6m7A1paCRD8ldECUdrQHpzEzlhAcK9WCCs5+alr
0zZ96s2tzyZMLpBHapt9UMU3YFwowitcgVly/5hE8iMUqk9pLMFwxegX09Z/eyAiht/cj+w+i873
9UThU/OCKFIEouxEIDyUFh+U1/HIn3EecrJx4wD5CDOioVaXTMVtMBUJPFSImvgGwJFZ8WQdjGzB
X9P9KE/oDAnpONCcjkEN67fV7uxPmIMidwYi9F/PVBquxPA7xzJs/l9UxBFU6RbshBouZjgJKDuc
aMAQHejh9FvHVQwRElF8aHPmfmGrtyMOBA/J2I/VW9UKu5wO0dy6Jmj9DtKQfSSzJB7HvhtdBS/k
wtKz8Vwf28A/4+gizV6IJvwoFvolAqwubPnVx4XLFVm+yXoJn1dCKjaJZzVTOkRtOiN+cXSFNOkU
0KBLM7C0Ef2EPqRLVHfaoIyLHNEKdF8JiO0BQdR5Co8vPRRbiBoKkqypCIwkYQiOMOFIwCoNDZnS
CEZNPyypjjQaqgYFh5CHRbdhBTqEnP1sQhsewuDlFmLIoyIjp+5a9MYCbSBPRCxEWdWL7grxC+l4
DXgtz3pN+qAwrHEO7l3kftBG9oltyT1JJJpYSPXFy8F1Vv6sDTC55157+Y9OTmhOIr0mGyNaqSgC
yq+ZMT4yn7XDyO2JtxevIlyp4ltR8xzkOiKYpfr1MQVdW4tkgjFenTssSkXmPP0t+Sl2VBs2Pxp5
2vcLZYIVNA9G6WjdfV7nGyga5hfErXcUX7GREJNSLURqh980AhLGf8rUIdms+IYdChNRmgg03n09
6QnZfhW3koHBkP1ORlgefB4vMiVIcYzDCnx1JEz0yd3qOahKnAAhX1K+EJoOBfgj9+iBhudmbu9u
eWlpL3OKmJ0Fb0FLGmUIaMyhBy4FZbn1Hc5lH5IVELrT5BK2yIQKEgjhjEmuHf0b7iZ0HoT/vMrg
2bhSxa0KjEcgWVcKiz9UAyQgfliYCxRhqtudhuU5zoLvZnHT66So8nFMwM3AMELGHrYekU9Jr4Zn
p58l1C4b6I23jvj0vlNob1NcOyFhUIA9/e5Yr09nGfyFVohvjSEkegzBMNT2SZdqHe+0L/egFmKD
ymXo5EAiyPMCxEz8RhkTYpFCKQXlYmZFadOr5Zik08UAqjK1GJta/oS76aQBMMWEUvTAH3zi511N
FYV1VhAfX/j2GF0PD/lZypXy8lim86GQo3YyPC96Goh7MSdCii0I5tBRUGi/rXM13Vl/5BYBvFbM
t5M5kLpkZ0pQQbBSi70rFnnoY3LWjWtl8fzo53bX3xEasuT79/JJF2hgdym6wS3HxBw7BNUlHEiz
C+u4x6uQD+QWNQWfFTfx/Z1FJc61Cx/zXuLfn5YM1ere6jdGrVWH4iPIbsW52MRSbB3/lkKfhEwR
iKkRRDpnXi/iv/Cjk9q66tWAI1NNGHJCBsFuHTVzWSuonH8vYAj65klUYfVOQSA0MfVtiATdizQd
VZ7Ryo5SD0zcPd00xML5lPxV7Udkn5cBcHm8Z/+I8PPRzR8w6ekcykh+ecUHvPe+mXnHpFZzaAhJ
i8GkwCTBR7obUNKWvy9BQm3wsarM9Pd/8OVmjbntVOgw1OHovdol8SViZbJM8fZ5o5cugurKq8+f
7tpyGwKrWwPda9QLjEahjp+XLC9H/h8lrBEDzJnhjsjt7jmVuDrEjG9zahgGosZZqDKcp+U5dI1d
Htlzly+Qk02U+mTt0Et4K+r7SbcJMx2KOQGOcKt5Di5DigFg2ugpjaSbyGiA1EoludBhsutC9WAJ
RJLa5Za9YNCVEcWGeHGyOkQE0PpjYUPnowsDqoQnEmmqdVGvm3EU6UfqzVtHEmOzaIMsk6DNGQjk
1ROhYyI166pEiGvLqIPSZXjeKoBtYXn+Zv2n4y39XQkNrD4nmgLS/kAcFf6Jt9oxoDGEFcFppHeq
+11VwEu1AwXSVkkBJk5ahTg0NCzM3ytEGxXoBX4XIZTDSKOUqy0NyvI1d36IEC8LU+FmEoV2+c3T
BUXf0mEIm8QGLLPg3f51kBj99rvycXjsE0JF5LHOP5QyAhRUd0Hv5zTVbrBNudg6FB6DOqBmEi4Q
7w9f8FBD/2A8bnkUBKDWAKjzs8CofalIiho0kx4i9vRZngQBCykbgXwqi8cPDeSBGqdHdRwpwzxU
voYDCTbFA+7vVqE0m2dWTxSNNVpFOqDx7xh9hcfnK7Vx1G71qrfDe/Oc7i/XJY/MP7v8nTG0/l3l
Z1vtLsdzg64qgZ++rqbo4dZ88oLf5o9QYJm+wQxu4sc26VB+XnXWQBlCpWgLmsWYV0eDFUTOwFjZ
C9Sf+bCf/klpS1baQX/0n9MNuCI2yEv8QJP2qCkUvMEimEBgXALI97MTM/wO8/7gn8AV5l4bFSh9
fu5kwyKxn4kZEfdI+OZ/A2lejX+VEtou9Ftwktksq0M8fnQftD4q/i/mWSrydPJudI51cN201gFe
O05daHzMa7oanvUJu0swRc6NXYQRLbjWCDMDr84X1ZaTrKZlAP9a4G02PUl4S+L9sBMJZL5zJ1/G
A6Eat3RDj29d331mG01/6NIxh3hSrrh6rdXUvhMcyQXLl9zIMs3ki+6J8S8C/+S1RqcmmhGuYBKm
EOpuqLhwYcyHb1fZ150b0GYuVGqWlLIwu7bUvHGAB+aw7F+w8ZBsiufCFBifWvQp4u8SlLweDIvP
F8Thpfj/xhsJdKDjntzc7jDagxmeLZN0M9Toj25Ca7+p8H9fiFA5buuEWLubnJdqDk7J4Rxb+o7M
NyTRy84Xei3iTb/q2cwkyPocjWy4UuVfFDYOq92dHZoJMW7rjJ70kqT9aV1k053F/WfUrdoxizuO
McMIWbJwnc/s4k1QMjOUKVkmNfyBenCxjYpcCLAhoF1GH2Cu0l13BASvI05YSxII5xIJ/xLor3lq
fHgG8JGaoVnV8xYYMSt46AyzPLwKusUhx7G9Oi2JTdbXsLXuaEVOgsxEz3Fw7RnR7ojPK6pyMuFe
1a0ADLDju6OVr9l4xTu6otwqRRo/TcKYJnE1SC4wNnVvhrp7yd2e1WbAWezEhV/VvDscrJwdEmDe
1S94DXoRth8rEwcjqm/Jnr6ZslLHLcj66oS8e7Q3COfOcifTmfYeVAKyeKHYgYoM5YxQQdw/1o65
NP5uCS12GRI+KX2KwTC0XGZI7zln8ryLDuqLunQeyb2UGcTY8LOz+XB8IEtFzkg9XTWLEHa0dL9R
exNXwHYlrfmEmW7/MMm3+Xu3/LaSnGioZ6+g1Cvc8nOBo1ymhVeuyXznBlR7szgdxNI4AFVzfNQ4
19nE9cFE37zUe0NCEN8eYoPYCrrEhZfJwL5zRg1bfd8UfhJgs1/TR8AdXPV2whYInfKoZGZJUsyS
X8zkOJm30QGrR7GMT7/mXJf8wR0Bhd2LgcTWzzvGSUXMj9LJbqV3s1FgLVoB2JycBvjZSC2qrqKZ
lxljWnsDWa2D4QZ4w9ATrqlPnhKKUpyF3R8A/DLjIlP/iqqw6h0FcMcL6UjKYWqmOiSBxbYbMEqW
vJtuSMKef8JuOVPyf3xTI+bN9WiBrvEuP0cu4K8cvuqIlVd0wburnVaCQ1+SU21gQCavoKIJ9UZ3
kgMR7OJZ/pVcsfMiVagnV9U8xzhswWJrSK+aR5o605tB/BF/USw1J5HIZwXxU4ofEyBmS60i9bsX
cUsk8wAobs/EA7oxUmJIo9pmu7dmwjz/gCW8pzqw764uMBBIpzO4nBw8HH/kHoVBlrxql4MMfMyQ
Iw0bHz3LttjQiqROgHeKxbgCt/TKNKUEuWasqkeM4XDWSY3hHOfsZWwCp0WXRoXrcxe/JOWcbofU
oBo/+mC39kVkqBrGPTyw0s5OuZGyBwdBnO/m4HyqkZQ71cLPDofaLFo/slquOtd4LF4d0kEcD0Db
Fi1rvaRNF+57NQaNI45MPJMm7i3jml/EPRabnVFfqKgZhei9aIH3zlwSrLiOhbRfKZDDnmUZtaRz
bkcHvnyfTz3h2XXFJDeIrudB0P9mErgKubkUyn3LGEXQyPPC97InTBlU/J/7zgrb7vtggsLKJmEy
vPlQ/2GRvy26Ibscsan3NaX+TUR02BUOLoIAiiNGAEU0C5cqeTH+zARcxewzKCje9FTPdK7I3GNV
O7ejbcxC+QvMrE+ADraZ6aaY8x2XjhqKCmkyb68Y+DjSzM7zoHLhYsnLa0SnigNTLsD8TutVmKiH
U1Q8d1l5wB2XiCbm386+Za319E16oBgRh6T8YWHJ+MSrLm2jpjNl2qSyYQcl7Cz+fI3yDxfe0lOo
TwdB4yVKwMElGZx1vrQ24jeiygCG4qAW/u6AnYFVALud75vm1faRgY/mfeubqgiHKShaavKoPx77
bYZDvqLHmHTJOv8/IvTUu/YcFYLu7FoT7y4o9y7ENE1cPufF90ckWiti65rUUMf1bt26iAuo7FEz
gLpcLCGK2Ohf+eiaeo3NuGrpr46DVqug9n0CnoVnW391DQzBx6KXJBad6ozX/iifIgtxFDk6MfNa
Iib1T5yHpIcxTF8QsTSjSAVj2smKEGc1XgR1OPo7dLkX1Nrci+/RB9i2R/xU91UINUBUs1qSVdw4
EKaf/qscraHdGqrAB0ywnCv/u5vblaZ9xxIouPK5jasyPTigXf44OE2ZBauVI7MZiJa2IetGD7PF
gWDWV8fAURmEUFD4wBhOr31Ap/0gw4taf3x6XJFF2iPJu0DIkK7chbrjdbN+AtPgSYlGinNIJSGP
Tf3Tq96KMx6Ml1AZvJTzlSD4Xor98KVyw1uNUfyESXaR++0BjW7Ai2uaEzyNP7DwsYd77Lteq3x1
QQOvEP5Qsf/Rb9KL5IYasMEYPnK/lufL3bto9nLseCejbfhOfAvz/gyvKYO3ob+cFsNVrqfw+41O
ERhINXo00L9AmZCGCwrDExuDqPne53kwjgfhmEa0piR2l+63/5xWZ/hHYO2oyu8X8US0yTtYcwNY
cSQXTYVR9wCEdbGNlO6LgFSSGcEPliTxq4TASUmqggC4lmp2XqIM8R2w/YUerogw69w5//vdK+qp
S/QikMwN5FSJM9bYxewyiDZjDdvgi+/6K1UJvX13vZusmp5OttG2wBvWNoz0UzFBbKgB9deId1Cw
IP39NvRtoEccKMqDhSiAgI/0/Aifmsi2pFPxt6B0GvBMAy0egVWqaDtJIbR+ePGJmAvNiNdUvGzl
XRRvIFVouBd53fM58Qowj+h9GHyljmLujUqMLMVjUgTDfARyZxMq/C10Lju1B0md9TX+Z1yS7AaB
QvCmjg406RZ/lCNYsXhKmamXK/ZKTN+/SUnhg3rl1laJEYmwk4Wbf03OxJS2J86owbYxeipBBoHZ
Kmt9MzLepi7hKWxOHOTjXjpuctjgung7sfZM2H3dCGe0/K7WZb2viTWJv91Z3HFDyDJ+ySPCOOZx
4RJKvksLcPJYDEe/F3KqD/+k2ZUtGEhZRxoQGn7LHVtAQW5U98oUE77hmwBPPW992xSP+BzOnVb4
mbDI/SjJzEUKsjFm96EPvMeA2Sgd0knlOXM1JBMDPMxQVZka2gGfMZccIekrTv/tTynyCSCpjJkb
jAnKWjV1VhIIwqlqS5lhT529PQCPRqeIExTHXh02oL5KHMnU8R1DzKrJRUghxOPbeHWxKWEuE5q/
nSdUf8RBYsrkFzaYCS4mkuBPhVwHO/51pGm7B2ZDZpGkObPkLDBJkNGR5uaK06f56batvN2bTVn+
bb5Ab4rK0oxq/4UsZc1zci7c+tlt7S11SjWXjFeKSgkY+JyRUA/3ZSzvTWgYGMiELVi+lAQIOwJB
ccRax6WemxduokTM3ekditmGHEOskmiFt7FsDKJkl/GEuU/z0BuVuD2CAAi9lKkTIXtuLSzcyDtc
Z/EdCU62E55P4Jo/BK52BCjCiPRprX29wFUREDhTvFzC37MPnO1yT6QiytexwfHLualI+WQ9WJj1
dWFID7aG4TXA3yNh0IhiYvsRW6ijQaaDEnpWuj8GX4Z04iAuqMZO69xdQmPOKmoE5aohXG4P2iYG
EUU9zd2FOr99RRc6tzRe4IIlyGLYff/NnSeE6zL0SeHGMoWpUlRvWoy5fe3GW25JIUL8x5TGd4cu
JyuKaOFEjOXOSR9WEQI+6K5UIK7zoMor937p0EuizmS5oPZKAD45GXHGpzcC3BCHo/+iLTKqkwVo
rwsxvfQV8/2Puw3F9NIwIagkKbqzoVft+0Dmxe5PSjF+ozC13HUqc1HSAL4It1AYPhbgk3vpD7OO
sXu4OFCU7RBYT3m1PmC035FIDBRB/VkXLZmAtEBzuVIT6FdIl9FJaaQ5AaxFwmJ0LxuumRKOki0A
sHz4HN7laqAWjr6Ibd6ua5fL+QmLI8/4p4HzfQo57o2a+orgioRuwHJzKBwVjNB8p/pUvplfVJMn
//bx1bCKAsXmFXMf6du9LCS2B/fko4L2dBPEZu/Aq12XcySjEwv1arQC1Tx6ox76PrF6sF6wzIq6
mMeZncbtNIafaj9Dtu114CSB/iGhR/Fc/4I5XpwAUDOkEzfBSZmujDgrj9BTQO8iTTnKPpcI6lRm
TMqlyH2y0S55Ebv1t6iO5thana/Rz7SGSXVcBmazTcccpp9iJGYhUiOd2kvw6F+qdx4RO1JIwVEJ
G702eHDTd4GrhyG9qGCGrPBcE+Lx+9FF1zRRxmGO764KaEJRZClM0OnxpKW39FwXhWjesBHoegzq
xL1Fbkc8WpHD9Q8R6hee8iLkf5iBEQs9Tjfgqn0WxAFNYyT9R0LKCqqgIjGfrecDBrI6tG/k1lIJ
WlKtEZHx3+RwEGEvW2St9frzGImJFzGXdAIDdI0w25OJQeUtdK7fm22USnQqEE07oVQdFkC94Di6
toPnfrvrA4bDXUChKwEy7MCLCoo9KXeDSInF8Ax4SoKcL/1PYlyY8pq/QuMUdq7g418WEG/2WTe6
/Tl5InUFeIB5Ax9tML+Sepry69sq6sQzgc4rrtxylxR0+aqav1lngHu2l+SelhrYSTRYSZsTMJP0
VjynA8bhWqDOTZLQHgmiqxKw9V+33BXrmWfjgv3z9LklqyviJs+fOMYGViUFYF3WSE9E9QHoI50Q
ZYm0DrSiu4Udt/Bh04eLGdySHJJGolqSjdI9aIGYzHmPNF0NNQpyZGOkmknkCvFLJo3EuPYjwVwp
ORPlc2jt/i5Ffcys7q9u1oAhNPSqjxaHnWcSfWK2+588+UD9nRaLl1e7uENiZY7sujMoh5m4LK31
tEU/Lj5DGDR/ljiJhTB0hKYFHw4CdJ6Q2AnuacZtPJDjH3msXV0WIFyjOXrJtolmSNABVMEaTuxd
Yy1Hj/kGsJ/yadwArhRUiQsptWZeVtf2dEVdSUIG2ZBJbOsat9G46AhjQ2bv6ZV1nKNs6LnfoRP4
3xb0IBKRE3tkxIkoFp+iNJOV3S34XOxef2csKii1yV4MYujq/5bZwrOr94pcZ2pn38gT779QJ56N
3qv7XrPi4vzYnTn9EzBkwjUZr1oqX3CrOjmPqXE3TCPdWH1PHkTNrVzz97F3FPYzmLRECNTuC9M8
QeSdnUajb5bMC5pHQNf70CVouBXXIUcDciLbN1dnlbyGyHWaIuko6KMcC22LujlS3SVRoo2ibkRX
jevmttEX5o1NxEndMzuy9xW6kwxGyasu5oCgPNyNaq7jDw+2b5TVl+t50T7zPFy+QXx0f4Ry/4/I
3QgBZWHavrqwDZOrgY1NO50F8BDhvNeFH/dPpmHKTekxpUn5pMdtIKHS/Yodh/s62scg/2XD5fmp
4ff8fbfcx81OpaF5SjT/jQzIjuqR7Wxdr8kjIR9q23q6mT5fdrgZ0a9xJ//CeHEvZsGfBYExL0r5
xSvxOyhw+8/4x5detCigACpwfkR7mErMBkgRjyXzLoh7ddUR6vSf+HASsqQafuz4lGJ2Z/rkIJV8
GkG5Wm2JdxfrCVw91jLE4TkEwdL86fBiJlPy+DvuG+cTEb0KSU4jFtzSrgzA29tqFK/V8T71ovzq
VwDCKlgPe/tLn/iVo95DoIH8g58pTsqJWUlSAZMwQuiEm6/zPbjp7q4tSLTcHsg+0ZX5fksYVRVC
JEc9UkA26R3Q1fMMdVbbi9mbSXFw7FW8HDskv9xIluQWnUy5FrbGPjLQBeZhd8cdYgxBjmR2dXDQ
QD8FYonoaSxv3EN3nxXkToX6Pbg68k7hMmtpRwIk5+BHg7Xs67lsRSzcg2UN/MOWV0EBxas06DYQ
yH5337wHfiliTu+I+5Iklz/JCeqIa4LgTfioAIzsynWXhAWieHzRDYsYGP2vyE2kZg56i/3/nMt2
tT+YS439N0pTNK9NbNCz5jPg3MmlRRIe9+idQ9yAX+TPr/cCgXZ1vCtWchv4UPwBIv/VsthN6N0f
JFRBWV5oN5+2FecfU+Kbd46FUIgMLG5MQ6IYHtJC6RfWtmALeie733Nwrn/WKtuxD5xmUdTESTvk
0SjGbEe6YTuBf9pDXCIA3LMM2IFtVXObbTyo/XOz0VsZ7LYd1ubcFNUJ1gTboOwvCbNHkiEMSOAg
eKo9uCZfc3gf0xRdbJgxWftQnuFBI0Pd71aSRCB+6j6IHI5OnhUHltYcZClvqTAW/NPz1uyR2hE2
HuOUG58F0G9q/wjgKIvQyLEbGw7YnJ6UP5j3Ai2lLiWtwti3dp1CUdC4SGrOznBDOh05C+wEe4/E
Hv49GsaywWjAU6HEYG1h+Cwej0/G2F0IQrN8QHGbAflZFGFgO+rxHZt0vfRx91SFDwLVzJaG1mAv
TR+mTQ16qegXz2JCN8rRK9TW9suq+mOsVEwq0LSNWSiZI8WclPdKHh1muLQV5snDRgaEbNopUxv0
Xjrdf11Fxv9rLjGH7KjKw8lHECbYygAtNOuKqraebS0OrCL+Ol+dqRjOkOhRt9LouzasR01g3Pt4
4olegXTPNnzV8GvO5telL7pyKTICqCZ13rkSSeYR71LcWV0NpYqrCaMwlTdxD6IEMbAhYxHsMA8H
ZXU/NyA4E2u7WIP7pSG9LmvZzoYpvgUau/2CG9RH2C9szJeQKtZe2cqay0U0us6uGIfij++3w8Gr
6dxZ9Vj9sNkBP+ocx5ZiocR/xysZDFUvdT+os7vIGBy+qnKThVqd0azsBkS2xziijnZs3JIZdTt0
5zlcRgYJ7XoRcFPElw5XsFJANsVXKkbe3DDhOMTr6m+JDsBjL7E0HLEdwx067nalL/rdpPhAXPXi
zvXU9BxDIU8lILrjQdl+0nMqrfAcv1ioZdJg9TxgfEGrma1p9bt0E2u4r+iVUJirG0ygQaHYDw4X
A8br+IIzbQ8JM3Z84Pi2iRBAhSyNGEXMzuI+d59jvswohb3xMqygSVTZzKbPf8KnNQZr90dfvKXq
6BzzFFU7BBhM/zYmJnxghQHtMm+fOG7H/Mi3eQBFgLuGc9V2EaiftnygakRSaj6EY0MKmCS2JgWD
JYHA0Ft4+CIo5t2RbZvbpiEPa6YAm140zrL6VWYmNbvQ67GbXI9AoKIayt8fgr9CkjGHJq+YEAw2
KnAfh9cjK7mC4pU0xsxVjUcDVfOLNuMTiyXOfxfKE3kkN4Mo5VWp1napkqEY2YO4Ew8I6NGM/ZkD
GnPVT6A1Po0Fiz+8Egl+35IsNldLyD814hdFh3OyUVswOmWyjkYVJDve9N8XIw88RCUaA+rLsu8e
E4kz9aCkThAwQUhnYX6yH4L/TywWD/8zzXNDa2Xvgq2ylgYVn2GjHjWoi6s6S8rn0oTDR892Kdf/
pn3zP7fbuIIRlT1yIr/sENWiYU+H8X7p2HvMWNV+eRy6iYYKXSqMpYbN+HLlK97H3MTuD5XBcHrZ
M9+EOA7cWhabNlE3CPksTZpxvjdV+p61e8dvYOaob4qGlPFF+R5fho4rHQwzSRw7kbPL/3GilO9j
Z8owmniTxFkz8zcmt/cYq9OYAZnhTrsFpe6eWEr4WP2actZNKL8gXUHVZWAzY8vK596CSpCIIPkX
PZd3QoKaofEIP2tbRDdZfRHJ6GgSdoiOIEWMABqapk2M+ad2IYotT1bNKi3S3/fEjWZYtAaiYhCs
3L5m6ioyf2S0t9FhlF2XF9Y6pwgy+1HG6i0CdeL0AMbob2eidMPrJ5NhKsYM2EbJJfNGtAeP8fkO
tGWueG37kq4wga/8Jg3/rWpaGBea2eFZh9MTxmb22fszKteQNLlvoK+QxSCaXKGmF9JCn6fQk/uS
G+H7cH+OaJzZtwEM0L337HHQG0/cvMdOcpTraP5VnaQ5C4a+0Y8eWmg7AkFkgP5DZXbz62KR5b53
XgnG5Q46XqG7a7pLSGH6TLX0yb66TYQ5RpzZKcxKbVlx3RvmanFOtJRZRamlWTgdHl9+GrChhb57
+OLVX5yreDC3AnRhhrdqUDxzvlbxjM7NvparlGiCGz0mxUlhfhK2yBo86n6xiwt90PByLRuXIyoA
7lXwEOk9r1ztC56xF++kPd0dDmojiggql10fQnva47KwrAZAGWqKllvPPVAJvD0+TJ7jNHFgaRQ4
1olGnpbsF6wq0YdeiNXT6p56duYCYACmFECpO7faCUgOq7AjaDSHv1cr98AsrXEn7MjgQ4DfOT82
VRkaGcH0fyfCq+TISFpFObrUPRNCU/awVHDKBPjXp3uYBe4pNwQBi19ApQtr6tqnFUgNuXvJrmiC
oaZFxxC+lUjmpysm0YbI5VwEYxYaoHOPkhNvwbTHjyJ1nGOMViHUWq12DFxDtpSQftrLRZN9ZMKM
0anUlRGfJJwFQ74Vdl+lP7sFfNmYqjJLRRnviHFkzLkYB9L77Zp5riQsbs49t/6cHR2HA19jppws
gmZTIjaT0UqeB53wfOfzDcQGQa9S8inCbTWN0zfmReyBvZYzp4b7UxggYvLmYILeeqzHo6ia5Jgj
Hdx9gcqWMW/JbqjmLVHPMWHQTZ6Pn24UjW4e7RPWbi4TkoOgCMU51JVQX5LSEyKovrCTlu6TL1n1
es0OdapjoGXp1D2NNWcZ0ygCor68VkOtRWvoR4syTJhcuV54gBpZILJhnOCyf9lRbmELzOaiNrAl
DfWTr+a09Kq7AfngrpbppuXjKpCjQWGi2qrLFIX/uc+4K/laKIdOChgI/jl5tWXZcuxH7G54aMb9
FV3gVZ+v1OZfzCan8YYkp4hpr8YVlp6S8yEYcjHuihyhfSOX7KX2mQPeGVFGVwr0Qu2zo49h2Hqd
I078WNjFLGCmcAUDHe3mcBOyk/C1tOfnr3u+Zm/YBwJEEMZjD7xBo1zoRw8Cy2CrM6OyfK7HhtCr
TiIpA/vJBTbstFh9Rm1U5ViISlZTgHe4a6jz+1iMcoVwC9XO+YtLObKup4ibSI7kwItK1oVrubHi
wW+vaguygWnPl5/hVHGOX5O514879cGmX1RIy1m1ziwjlyfwx/apfCPQ3M2paVcDxd0FlmUcHprO
2m3EGYLo7jKrDkIY+H0G62sW+F9HHuIMBjVGZMbk9TESwW35MDEgIlQuJLntnbfJ+h2lnK2HTpIy
vaml3E9UuvrK9qG+ltIv/x6+Z2p5lgReUjbE+23jYm1bsltF+/+IfieS8z8tx660KyDx1LYaEgjB
WQWWPYfKvTrbwC7+Qi0ySqs8eViVW/4FA4rF8x9pNn7x5gTCmrnIjkR+uJqImDIaQw28lD2ef+Td
hyVAFrA9H8uw2WPd5DalBg4ajcX8roC2STZagM92Nji1x9V1mRzkz+J8VGhxlkKVXAkzTQGZEPOw
x+0z8cn2Bpy+/H8PzhnBm47O0nXY4jdUNG1O4ckQPCCvfkXZrCUYCist0L5lZxVBtA3jN/sgx1Iq
uDz24Jn+coN+PgChUlWyYzTa4xxkEEA2tG8UfFlge+uHsoBeB6jYWtlL0ZME1vrhweibOrCs2jaw
NQI73B76MOkuRhq1dIfbZkKIa9FV/biIErZczE5zw2wjBBLlLKOe644AfnAeFB8x6JjfJBP6eHUW
SM6V0e7K9IMyS9tFOcsp77C6ct6wy3yQVP/ULgYjYvSYegyfVJ74uJMgOkXqQ+B0RTTsmk9q9OOs
HyemB5fccv3V6FUk50N30Sha4v26AiNOP8l5IGUEvm/3AB8Wsee1YZUZFRX5I++kz5TXy76n4hgK
owzaBq8R0/1eqkMrYlc2FlhRU9s8mLwRDldVRSu5kRrMLmh18oCj1Gd/pRHCNBedWlY+kxCkjUDQ
7J7xQW8z7LxGryMCVDUTlcL+xofKjvdEIALIM3fhp2r+pfDyGt6X/fckf6rg9q9dL9+oaixJoEFL
e+DoInW2jYzctOQyluTGMMtOKeI2j7ood+lCAMKbeQGhpdI44xG0puB7UT5wDqSiAcQTQBtQ1Kxb
8rp76nKFpycJaHioHGdl3aQYV98L+MLzLdQowJFUCFCXA+Js7M7z/91fYJc8+NYO+k1AAM8JYRN5
ttbmovBTE1hkVlayKy20JVG7CqwZVtLPASCnDMu4xv7GmvO3jb1BvOMnSngUgRGwvYT61TX64F2p
m79M5bppr/dAHvKGzV/l1Q8eaZP39KRw8Lo/dAQXXHu7XrtpeYH3XZfX+/08IekLMk0o5B112XRt
cuXJAa7RlOJTcA/upqJCECWR6PYr7JPeCwCBjLeB4gsWW+ueHba4xuKbiTbkpMFn+LCmMA6XmhjA
/t0DeyMBiXj09Ts9v2YIzWOXiQOD348MParDstqQeXLOZX5QKRCr3nuRm04sX0+3hf082SAIny4d
jwBi2gwDOt4RLzOntAYaUT9MJMlZcmovY1IX8hKWZ/0aGxRIGCBNXuvre5Y3Yt7HKJakc9M6bkmq
P2/lc3mYZDebHE34955/oH+2k2xiKhazHHieJ2oghfFWEam67nEOPJORBCxX/Ee8aap6JnPBl/UU
tkC5Bx1X//7fO8kNhSDCOvdYTbKTqeVvo9FwZC8zWDh8zdvBl2Pazd06joNAku3SS7Gn4HeyODwX
aCOlOgPOerGt/ipaTF7GpTqKm1UCgpKCPxifqcvAhsJpGibSNohL0BWI32zI7x/YI5Z+G8SvOy98
LhinzUosuYif+anyup6U7Mb3kp/tmkjOv+mmhAeUFCq+vrFmWwRvGpfDEC5JH210nmULSmVTD8CA
pXlc74bwzBE5dT44UPlR4AbGAE8bXX2pWF3aPXsNCInzvKMQtveoft2UVMiUVEDdfndaThxyqbER
7sKQ1vdMrNzG31yjYWkZCP5wRdaQvdTxGY7iuNuV8M9OqRZqoP80nK9Dpx7TarVIi6skKLa4VSVo
uYG+5Y9rR2xyFl3GtufRUvPal1BbDeR9r7C7BnIQ9qXSbdSJin4n8MBnW9eyOkRfCkRMeZYO3nRQ
5Oj0ps0BJpKuAqGAcJGB5ySMNVLT1iJk0i/0CWvpNGnTOxXEBc73spGf9MW1rcUqaqTTFMXY0ivO
/xWhyAIS1HWMZat5Rak/llqEnIw/qgkQOagXgou1UaVKvIbqL5vVSY0LMyL2EorLdZbvpssDZgLW
fVeuuLb2UxF70zJh8YHhyCcO8usk/1rLd2cWfRC+aFlkOVgTkEj2YJuukkuVQgPPCRW/BQOwwXze
SrOcSfglqkxbxLLGuCvBSexZLLW/T2K3Y6zIOXiPGpog1shbiYRrUXfSgauUkQNXhS7LepcWF+Zh
P13KhvwQ0tkXEbKEsSIp+tdhKem8PbgtzoCQQUEpe6NhbSJFwiwL1xUcudVG66Ve7JNVqERiSCjH
lMlfOjSzxQdcDmsLmU2AGfxopuoWzRhTvsKdSv2+2ez9+Lr/j5NlQJShwrRLkGYO3zQpRxnDCvzB
KbJ2QpnO1xooXJ/aWH+letB2cjWgOlCxnl0HImeF6pZ19UNw004ZLAKzDGdW/Ry4evtjyoCy0cfa
CCbyqLHP1zq6tGAYR+TFz6IGvQL6e5rBISNVjR9qCLW21DFphWx6cJdasLlQd9pvT6brjiIluAEi
KpdQ/QZwAm7LL74j0u7JfRcbd3wRnjYEfnWqmUNHBEyaUEx/G7M2RtlK708SGYDb1wQqboCuxN03
4WRkK6iEKtAbFD33e3HjkDvrRIav9GQzT0w6HFeU7WcxoCl0fkRHxV8fYjm1I5OKL3CQxdr5D0aQ
2OvnQ8406iwsSUp0eDYDYqvYX/eWF0awxvJwjwNooCXlK9tMtPRxkoCaXnKVjA27/bcsXmpjVUy/
tD9c6uljNA9E7xw+sDrTR4Q/wZO8aRvF7D7eKfZ2iLJWx0s8Su+sXBpHhv+4177v0fqprv/+k+Va
zhGPUNFLrsTPwAIJ4ReYwqQ6jYS+Kgnvt0z/LxBCz0ojtuUMPhhva0AOc2hSqfQ9PYQ3WEbEy0SU
06nbY14Fzyz/94rsX2XCFecAOqPOiB7woiX/fgX89pNM4HCgrDzThLTrO5nFbvLfa1UE5H0431mk
UtLv4hKsXegkYgQTdufuLIHdMcwjNzQ1cwfox9AzDly/XxKHr2GNnkfSDq3oOmtImFw0mV6ntrYI
fItV81KGFGlo64yjtpy8G0787pDY1R4itDsZNDioleluAZ1H8tJtFBkBr4wZB8KEh7W4C/Q71A3q
g1NeQFPLf57zilYo/SlZPdwrxQ6BAsuY25m4mtqlVpjDZLQq4SfNUZFEzqooGeVIx6vhJivXgB8s
svD5AuPpJGeXR4ReB3QlOUr57We1Z3o6JgDN1HODWDsj7Dozxny44KcCSinaYH29oxnrNm9sGedI
gl4lMagQgIXw+3btzpafqWLsiA6VNTYbdO7m0gjDxEII1TRxSq8XK7JRPXjY1Jpu81PiD/cju9aH
wEkyJOR9KE2SjmnhEXUCtV8RI1Z6Dk1mt/1TrPBjqksPT9HBTUjEjdrO5amolGrQAOuOVHQC+3Mq
Z0wrtHIq+40IE+/ZYpFXah2SpCvOa0iwKSb1ucmtuQx4IgMRG5jj5wz0iAwTI5XFusEduqvzGQqQ
hv9QKPPQkgeq/SMJidd8jSOor/OkfKFS/uCoGVA4dRSMWZ0hqGYAF1GkFRDTYZEWOez3xE6TtTnm
kAJ1ROy2AXgPpG1U5BkvuBTb9p77enYkqxvNx3ua2fIuykHnoBsXJC+xs6XC6ojWtKxtn4sxx7NU
F+zzJRrr5hCFZ22sbwXtccTJKlhVcq6lE1+o9h7s+POAwwZq7DBKTpPdkMa2Jbspj5iFSJXTbxOm
jezSZKWPZ+TX9cflccKtsOsc6UKpJ8Xpgw9ReBd1xVHJUouP4w9Je96YeBu0cKCEfalwh83efjCz
BRtM0RX1stdknc6Kd+KmSTtQFrSD0eP+4rURqxIHopqJdpgvsBFRL+W9C2IQ7YARs154drl2FMvB
rdnV63b43H0DbyuZ1T17X/dUHWoJki3y/S8wv+Dc0v+d8+2w3mbbdiko6HCHV4EzWZdd68lZy1yV
aZa7jD/5HaV+EkGl3j4kUgES+WA/3LzwQA988ep/bpzVslH6x7rNH8JZpX8NQSswwTH+y6RmkZ7j
N5xbuCR84syTdjS+egJCxMjrggEgse9/jOVkfD6A5H8thfoMy6jYBtr8OgaxJUoZ2Er3ql0KfQCS
Rz/pnsUOg0f6vl1OyiftI4r2aQfcYg9EVYTIsBtOpgAJdcTTr0rNKmFC+vX7XgTSEAi/0uqhDB2c
GomTFWyvApWQKI+u35NXLBFLuXqa4ut8prPzP0NdkH+wZDWyGylEkw4rL7SOgYhhpbMm9OObmnar
j2CTcdOdYGebLo2ETKDkvXJtNnqJ3m2I7Vm3Pdgb9p2rHgox+zh74BjztEurc/c6aJfMdm0ekLZK
MPdZ1A+j+6llBuGdlBAPM1F8s7ydPImYg3BUBdrBx+7k+wGEB6nd6Wq0a/Z4ZMUljPcU3E3L9NRb
pMJ51u9TEGVyfnBvoYHLFkGzjh58iH30mJV/22QC4M0lAPcTZgW4m+s1BFJKbfuwHJVBNiXEG4j/
jY5pp13ZeNiN1A8YAx8e7sPkbVOK7EazU23pxqbioEpUU0rQVeJLMkuUwySPxzvZ8emna3MSKzOP
apkPBBxXBAIag8LHEifQojEKXzuZ9wdpd7WT56bEltOPlCoBmJZVkri0vXiwHDXsPM7+NE5xOIDa
HOl9mN+6qFt1thWmeu0Zwa+Puy9V1AcZDkGYGDpUnY61y/UsqDOsVMp1OE9qfWURJSgO2n1Oj4MP
p6HQRQALKaf5ek5FU+a+j3i0HyEuW5GEW6ObxIZggxuVrWSZXw5myRlBgIN80X9cp562nvONTJSZ
NdqJZl83ZBlTlEr2zeaXCwjBX9z85k1FwpVjJCbEjfNnuWtYuCzAR4k/ePai/RQVFQD1GRy5yr/c
TLGURIPmdFNkaKwE2VWLYByIxRRgFPzJ3zimjAeD+ql7mTPH866ghGiLtQLAZyvSx2PxpHqh5qO1
b40/5mccfux5oNN8mXaNl4nIveFdj9tlRYJKjZLKkqHjhzaUqOvKCKgCnJeQdmG7esidKf6obaRj
gUKKb6u58u7H0P6WyTtMx1azyrmZyOJzAS5MdtkvK4hqncp0Jm483vLaayDVUoYA5LyBNbOaSMA+
WSoQaL1yQNAKeVqaCu2hOv0iZ403sPTw30Awbw2nQpXOcOnKwuKgEz3xdtyjydvOX63/+ar/mzdT
2pgvVJYj+tT9bl0nL7CaVYOOvDIuATgjjIDUC8SvAA8juBcGi/7XQLz96lblRgBjKuhuyDpkxX73
7EJr5TjzClB02jH2w+Slo7R+fh56qQ/w54ILmnE5gruxIQMYxcgXNb5qGDqmC0qxJonbPvRi3k1o
f8kj119bHJzf+25IL6ZNdltz+IHuwmFJTy6rgFNZ6unoWjJgC3/SqDGOb0dGwJ/6FxYa38gFUCPF
9ku5RpUzDKNEZrSCf0phO4BwHTI3l7UXoHy/uJUupXu8G53C0GiYSOU6baubjEJTJ+UypDgzAfYN
F/cX7nunk25UqUDR864Gh7t0uNJJu1S0S3+fGmUSyejjd1xAXaSQDBKVPg/WMpytJinB9C55O1AI
UtXoXEHA/Ev6A72qznGXV/Vkjqiu20v5cqlsLiApVzNyUUTcUARx6rWQbJIk/M5LSpa1eRic4rVV
OwJyjy+cnNCUfCnjMUDFK7owZOpUhXIO3rknNu5Sqd70QtlSPAcSwr8gIkGQmFo2Sv72dxbqSTxs
zz3bVwG8sdp/8pJa21t8+L6KkMjKZug3FQKu9wkOIkqGxfSHmdsOKec2rquDo2thKQrcXr/a9zYr
8h2v2N3zyNCdrs2MU7P/DL9xKjRDBu/xeZvahS1xdCWuO9WShqTno08Gah9c54Zcg06kvFF/M+dX
Xzb7TuBAlCzXPrJGeTvPmA3TRMJOPjZc2T7hSJBh+OEFfL6COTWd/WOuvo58ovOMMRrsE1VjzkgA
XBcSM7oc5e8LhfPud8S1M3ya3AVpvSZ7VvamdU/u5pvQpXUbF8ccRlddWoqo1lxPL1caQ93t3DHq
R02kiHEiahAzORRUttKD7htOOj0InYypIpzBpUdqGZhI+0hyoVSSQQwszNp9AAzW9/j9jtovM1Sf
r5Y+MvoFRenDmEoh2ulr4j4XBB2ngUuBRwbXtGBPQXycGmieUUUtc0d4Ufplt3uoUt+icSWgZTDB
SDPD4mdwtIvRYkhh6UkBWlzZE1HdaRWUTeOJt/KXE2YZjyQwQtpJJvKdNjWqLWblbGpf7PIDOFBp
P/Txdc1r8PBeVTt1kco/a0vkNtYn9hSry5Ff5yU6+/rz9+uUSiBvx01OaotUDDzk81NAQVsasg3Y
C6qeb+vZjjmIXMu/KhkFehRzTGGDyEN7gLU0QXidjOaA2m/6VaX6oU9uR0p7S/h2XTQ9D9d6zJML
erowfqMj0QYyrNhFCffnCaOJqpKZeQwLMd2XzwvYMFxmhB45SKbh1A/018PuGeTyIUAwiLB1W+UH
GSACxXCtWzTm/pI+DWdAZ7uzIDEz5oC2rVE+1QxwbN4OxOIGSt2VjyiES3SWrMm0RnCt4iUa13n1
29lswQluk+TOXTTqkSXRCs9A2H3B/3DVgEGl29ihjalkkGyRMOeBBcv3T/zzvyMEoDtb+IJerUz4
QU8lBGf4Y38dPsHJeCFjhmLHQSRitGAvSQUTD8g7fjY2gcGTCB2isuyovNZ6RC8L7JGzxtAnoQA6
djmivvRDYopJ9pjyqZVz/cQpbL0J6mMPL5bZ8x4xWvccIYdRiF7v1pc59lJEdU1xX286IydIGW+i
gIUpora+DUJ2nIJ/Q/xuxe4xI7HX3XnB8x1bCdCLGujq9o4vCDtcjrYo/4pBch+aE1HjF/ml4E/Z
F3d4SL2jFC5CEPSyYF69Pfb8AtXXlQlHnMmXqzo6kEQpncLK9Yapp77rOoV5OeKl3VD5ZgkP7URT
J3+fdaZhFKp0yoOJY2DqzZcAHdxJXXJ+Z3rWpKBqMbDCTfBbllQfddv8fUCpMgb2QWb50FA4NcKS
uqokWQtAGJ9PPb/qPyx/7HORVt4M89EGvLu/oA41+omQeZVlyRsOAcL7k8AGkAgtcj6RLjRvB6kk
d/zMJ3XduWTeD9wFCJ5S5t9N7BJ2sDH7S2wt2oDBK9Z6fDBdsQOPU6XIJEWKpH6gvrZz2FXR09da
6pZOmm2xkDZEUYbuUpCje3LjTiaBu5VQa+47bAWtADIMXzEkfaZdoir198t2u6Ed38DYGBRwAGpu
aFK/EIci5i1Hx2IntfXBnn9UL/eXWO2nMUdB0Y60WOAXn4k+OsUGqvP5Hvf0kS36ug5lYxsp6LRa
8IwkyRveMJnHy0wKBhvdXiG/E2fjSvTfcdTeHIkm9izGMeFlXW09q9Agbxy2XsQ/AHTxS/9Fa9X2
uFpUUwjFYn5AXZEjRElZm7TpK4VcPM1KpJUUAbqc3h4t/mP6G6AodW1OFbpELCD6NJWKbrYCnINQ
vPcMZcN3O/DobNr6OO/jBrDg+kUCepdcniYk0EmRWgxgQbz/eA5d5xrJggK5D4ertuU54pgNGUcm
pl+EnXjM3Wd7gOE0qrulDPGKd7h59oiQyVMLc1PtqekyK0XUJXjybKWcBgOjhwNr2z5EB6r9HgjH
WYIKi4Lkt1VkA3du0nimy8WAxhU3b4DZ2dvDFx+sAinjmL/Ec6dGCK4HXcAga566NxrL6md+SrMl
gkwSHRVM+nSOrcKou5f9TuhfndEivl4M2wGpu7fJeYEOk5n4lTHwKhZu0XBMAL2FuR4+yzAVaI7N
kmJ8i/G5UIrlAU/kcj4HFTM6UeVgG6haYyZGUJ9XmMcyi2QNMZnrEOLWdujHyOQV2gUUwjTIbq0I
ZqVoWAapvjmxyUxHLKi+8GXTxJy7CVU+sHNNkoXDQqCj9oec4rPXD+VKYTwFJxZrX8axgXKDC6ET
NT0sReWboGFr6PZj+8A0VUleCl0zWQpiPDZEgaDeBArp1xQ9cOaFTwvMJ0nOn+79QmkU0YCczQU2
HirHkTqJDzJwCFXSN/ICH1WPAFTuxEqmHKhsz4HNmGrfUIVpWY4FBIzkXqwoWfHnOWTM3KIIMC9x
PqfhHGrLxKPlpvPFkyxvyQ6tRjBmLIaCvl3j7VBxN3Ghk6GpoTmVOfHbvQ6SsrfIhSxNYgzfytGQ
RUzrstvyLTCu+Odm52oMho5M17zk0CxRqMoxcuLEDJPJYfzHfM65kleqarY+DFo8jmFUD5P81cDY
HU8POXetSZyQl8xVE0L0gugWZbyYu5+BA6l6diyA6NgJUffR0meTDkxm9ac+iU0p3iOT+uqIYsvl
Y2LT26d6FFPe4+2ZNk+WRfzB6q0THbFbjvpUG2SPqa+dNy7EORW8bosEbi/qH8q2DgM/9AuLQIwg
aubXeSsxKUhmHXZ30ohllZf48kGLncUZXZBiC2wk8f/UMkgUE0uOhVA8zIfhHx+MzwfqM70XfDDU
cyzIbSGUbqlRfOCHiJh1gWxinTGhmqwS1lJgbuc5j2kCYdY9CRq50Zn110vyzgCqg39so0CvZLLS
12QS5flGVsRWoERCZssk81P7GNRyD7RZkZ456/es4BvLxaGWB5C2K1DvON23j/oQ+vTq4SP0qB1F
LOlPMKm6PxBy7YEZ3YE4UFvO4TdI6TTT/psGI9GZ8SkTgTqW0Cz3xlbdOK/AQBxE7WOZmPT4SSjW
BN4i74Q0Az2PkAEBamx6NRBvtUTJgJmNtEHoHaN+ibsDB9LXs7hAuOBaRuS3Kys4Yjj2YoE63PGI
KpMUXuAPrKwbcU+AjxQkmxJw+gQwmykm6vNhu7a9VXlAwikMsWSqvwzViYpQgTj6UXgh3dxRnNiM
nKQw+bdW0p8DYZbvF9qZfEoZpZZNxyajGn4xDxIuqB+ffMSwNoiUFNT1GXu5F4EN3bKEKOE89x2y
tCpWoGDZGNXuK2lgtJizH1snqUGfHVIA9piUc0sXUsn/Xqhp8hraoxmu14ArOp1ha0VU12+BA+t/
8XPebZgX6N6uf7esU+zCGlMp6OecGDJ6jBQILu7zM84YRlYz9kKG5wedfCBUJQrL6O32PfM/0KM7
Xs6dLI0Hm9cT3vPTjB3qpqddPXy7fJ3nfX2i+8lYtLfBa9wOBDSOoAdU6rzR3vJOiko9btta1S3J
JW2z8atpDd5Wimp0SHIxBoR0rAYqIlOBFn2STlB4I7OUIS8UiFdBefWg9sakQSdD9PIDAxBqQZWc
hj2Q1dfnOnHP3sb8VqswUsaMRAjrjlA3emWaIqS5rHA3+r6piI6Q2FifIFuvzDdhfGqcRtT768k7
AQeesVZGQYWDBpwzxB26aPo+M7JdBjPJEqxohFGu/coLsS+C+sB7e1c6TFoR90fzPG6RVFAyWZix
TCn62BZao+OiGG11sri+TTHobGUoKVFmLAAeWx2E6nj95I4njSYBXcl9quAK2hQ/QIklnXFLRMyO
/qsL4U8lQ8yICf3Z9Zo/GWV4d/851G60sBRNUAy/A07kpFiQlEsDAcIjBEhOOtSCiibFphzGLCqk
RtF2qNlM2Z6gLicZINyUQOrANgJgPMrjk1GKTPgRLGuEd9N8du/z1YMKiGulCEsbTNhUqO5eevhV
9yvVAR9mmJcRUaaNlPICheqIa3RoNkjBUs1gOL+wHwUG1m1KoQNbgKTiDQh7of4sljAP2AYHPeaf
0zQ0SO1EIJ9TQE6x7FKkFdUiWFNYoYijFVlGTp4+AIyODeiANq7gS5j62ZuSnpSNEvjGlXZATd6C
l0iYEGd4taBwZ0yb3N8A6TarXAZkbqBOvGVxEtJIxy6HX8m/CcN2VrWDOaq0cIoHWCPBkFDHgx8Y
Vqp8Sh3KNBAGiDAD8H2Ix//+ofxaH0Jn+dJhGTDr29JxOe3gsCnG4sIC06lHNFhBXljqshr/NaQW
116QzObjtdT2QPRa0rELnPYqVNRKeCZlJK8pMTG4OU8c5gPRY5KBkaeoGQX4sQSNs1vg1tKL0bFS
a8L8dtRXJG6hlnaAS0HKV6Ct/EeupwF67xDzuJDa7PuYfFdx2ck1KCUL6zpYkF8VahRNdEwHDloD
a79H7sXo0R/cW1TEq9bQNFEh+EQtFchHlF+j33D85i83XY5WgSCm1KQgPFRx0xgiHOvpQhkBk5aU
Jq4jx0iemxGFVV3mntKhE0IFd7A0uoy80czsEYdPhxQv6GUNQeNdcK3CumlaJhPoh0Fn23eXDsyc
IegyZOdfGMpP3hCAdtd+QuA0ANu6sXBcd1nUyqHJxHfMrybz/YQGdI2YjNsILowGzUJBHTUGx81s
dKYaf8y1+jI/X7+0JiNT6VdN07tBap3oZqRDea+OfH7YxfBh8dwi0zO7BjHMVPztqe3Y8sF8+QQg
LpISwcnHHk9n1/s7e6LnHqFOW2AOBGEnjKcESbNs/ckffBK2tfrXEFr6ctNU/FJ3ytmW9Y7dj3yM
Y/nj3EbpJa8YYZ8/vpgx0gtkeUD3KJrx9IBsOCwYIJ5Tfgljftkw+/H9z9vKiHAzn58OqHsEt2KH
+Ya8RL6ZRHqLU3S7OX6ox5cKDC2ud9ESS5dOgikWL28bKlxuIDc14JHprzuoVtkYYNQ0VwEmeWgY
t2Tffm7CqVvok8IHCJIqC7aIR4eNmhcAfPL8J6I6DlLzcx81AyoViLNrP0w3ow+n7WfIASPyEnex
E0iNdnEWeOKwc0AHWWByXHeIJV92aIoLmKJxc2rnEhOw+QpEP9fUMnrz8jDvj1DrXsgC/Md80N4o
QqnLevYyJjsPndaM4rh+GFbrMWZ3G2h7fTaWJaRr82MoqeZSTIeRrYg+ZSPUx82AGJKPHTtRGtZz
w10CF2/Yo5jvSx3v2nTIY2axmQgzyG5gCRFxrxN7XCXhjgzkeyDEUfYrcIzltzd4VU6QI3LjWcX7
kJ3a52YLX0ocYmjFsz1w7GpE0LwNKXlBPly3JPjHTQkZO/amGxtKcufEHfTt8aOhrt2Gp2C5rEeO
Iswin5mxXS5T8WWeADd9BdaE+0zhk9xzVcnXZUP5EzxeQ3wOmRdiQhMmW6tqcmMNlQQNjw1QxZ7b
gzOfc1CKnX9F06o/92SSylvdN0/GwKTnkfLQM/MB3zgzehGGR+FZp7KxVxGLeMnQ4TckwuQGfSk1
03b83SDRGH5Vr55BbuwgEVWaP8SoItMxDRYDf7zLK4z7+PHCoFTsN5+IsAQqf5sjAHUgJblRTnSh
gS10uSKNp2hU2xkxjQ6kmW4NaUH1SqKyb4XyTmrmoL++DElr96ZlRoFOTn70Pn7DeNM27c4rXPGI
05WtX4P17EDrSCdjNDVOPA7bexrSxY5fuce1jlcKZboiiXcl/efpcMiCs80t0UnzF+Jw9M+ctdPP
JwkxHtyvfiuus9tm3gGttcR/jKPZXOcvc1ksD2DdaDgjh5KTFPp+s9xOeBsLjgpnTmn4nsp5eTyu
qwJIJbtf5QY9a/sPSkDTUT69qzorjrA0FWMlePpm7jvv5r+y7Vnw/mU55GbNYEEoidSqUNmODchx
iqAou8l+ymg8haYBx5ClC3ivL83NwCfFonA9pFrChHe3ihJLGy1tJnlBVTX6qfPwTjkxTA6SnsQL
DoJGumTrEc39iMSbh0FLSPkfybcz4VOIKe+a0PMGIb2FY63n5aQGtpz4jAg3tAk0ipsF1ooNHOBN
xpi7UBZ9kSlnhZvUySSLf7zsw3H7VLgWxpbJ+ezUgCso44Zei5uRIUv0GA3znxWVkkJEanOoBBeY
sAtuFY9nUSyg/PQ+RRZcX+29jrmvz1qOfygOCUoj3FdJtdxxWU2G2uOYn1iYMDDCpobVwyw6jz1J
p8YY6K66D1MhhudjRWpvmlpYBHhMVlge2tlm9wqkBEimwdgmJmyADA7NGS2RHhbUuWiqIBEA25PY
rkQcY0XA/L/iZkzunYLg24n+zlWKZ/l38Mory2qGXZ3PD5iuSCmeFc85Fp1ILw6ajos3bjQN6jeJ
D+t33PqzCpCtsxzcpwJBrp5EYyR+nL4QMlyAvusHic3/jdraQR/xPeYIRvmXKnvV6p0MBOQR/PuE
SCqhSZ0j4WktPYiLygBojNdh6LRCw5FQ4LtTHgh606fiLZZPB1ugMNRfF2/jooIE4Fw5ziAarj+H
i451uLFc3fNvvzHphQDSZChRqeHWrkq63VVYTNSuN/0t519Qs/Ern/97ZzUk9qsqGUBQOl+R8Dae
XxnGHPMr8NdljKourIDhNp0uLlpKIma0AIwlZuw3AK3IdYEPQFM8aSS+dtCmrUnIS5E8DvcG1t/J
MeEydBY3bpBGnAZJnuQ5ZCKbdX/5NY3rIAh+hsx9iay0aXoIa2201BLz7e7xL636HNVfs5OsGHAs
nS8QcHzooh4s487Yw4vN5VoBhvCDQuUqPyaEImkPgZsSCxilwN4+PYFPImBVhqF/nRS+kQL/ZoXt
34sRG5csz8a+jK4hyHU18kWhbT8kxqFn8vE0ot6W4QB3aVpsoEaC3xATqLEqtnWGc4F2Y3JIIAvD
u8DoaaUj/wRB2cuZjchpNCOM4DGOFRNctRhz9Zkt2WuHMaetfGa2YG9rJMcsqzrDTP7e+MxyIm1I
0SySpPJo5pjLlFh7ys5dacRLyFBqxjACEm3v53MRpJL1JBgfsLRp4XNrFk0KCYV7h39EKo4iYyrw
WsiN1dqb8JLAO18tjQWHIvKvh7TotRK8MPOAfY8F0KBIPFfbeaM+8ygr4BOMOonMX833THfQB55O
3q8AAazhJLO792sYI7mAU7ndfECgEAF6ktkjepjZQhKzfLfLyEQmO7LjH6oOpuUEy7fpY4DUE1T0
isaJspnZrLps4IxUGI5RwFvns+bBXEvIxeLy96/gMXwZC31aiSFV4vvKUoPn4E1lfSwmFLqwrIwe
CKE9dxSebwAehBCuXgjj5jkkUBYqhHSa97nraYULndplX3X7h+D/qG1LD6gK7zI+xoaHQtpXMOqf
WL3bJ3TFNwrByOO60ty5Uw8AEYcs75sAimhyD5Iy05g6js9SG67Pha1bV6IzBkpBf5Y+e4VjQFaM
ea6b2jA6jd4kNjPjKY7Svim+h1o0YNX08VpG55z709maDQFOIwhLZedcYi7NuOolT9Q+ASsSWYLs
RW83CV2Umukaz0km0Bjcc1pT07w2T8XcohJpPr5oEGU0kX0YXj6icfPHQL9kuB9uO8sHQBKyrpi+
g9z3VvO2U1NROBAeCVRMyVLMdBlxtx69JU5ySmognNkW+dAGhROjR/k3/pa76XtT6M/6nn2nPqyp
fOiauGoiOgUwua1DxjgktCLysPIIKpciQb5r+kIFDPFWuwLQ/FmVZacZnUp9jXHQS+UaVxKIlUcC
YiHTY+ggu/R6qJ02bvFCmDcNBdemo0Ygbt66Xa9YJaTgI6ecqOdsVv689lEWV73hYRAA4h637hRH
zMdJ8vCv/Wy7EdTpFwSoeTJPrHZPXP5ctvMcVp//rXl1MxOgLJvfudKDddp2UmgNvFkC4LFEno7v
hQMoO8kszh3t246Oc5m1Lj2WasD+Uq+iKf6rz5QnLuDBD3GnPVUjw95EkxjQXXu58Jzy+pVyZKRo
a/dlPrWAjB/n0dup8wbjnb/opkuOM+Ez3VrjL7vE5WlMU2Ch2iAnTIYVU3nkjUvK0JNdCADPzT7f
k9txGMW52AAFPU1kLKESKqeRCBdo8zqLRKS7OM1Lxbidri/eEWrrTZxziTzF5AWXs1G9wmhYOme0
bOePaCiyDuPyoKzQBWMgeyTeVeMdLEtvOHMKPaELYus4GKS9tPNSKehoq7vhdn/89HfgL6zCKJAT
Gz2T9vySRDQdtKW5Whv/zo9uDCkA8eOhJkvjMatrMETjGqa7pGxxES+PfnWtjEmrErNhrgiFBr6A
izApoZbK1aoOW1kG3q3R9A5YQAMm8vei9qm/jJA7/S5QtSWdKvQf13mROI2+D05QlwbAFRIMqN8e
rVySBB4zJcXkOdLgvA442yKs1ViPnmC0j7hkCo7FPS5zF5xrvBpCSTGnK55W8QlVpVvQkuT58a8N
wO/mCMgT7c20RNu+xxhn3jK0jL/90nl7MZ4RscOReoJN1iroi/z/fbSvuaVNlGOsf36oGhHdgX0h
dEek7GWXidMGPn1T9jRLo2R1DIEvMxCAvEdg1+MXBI4WDmTTqFqMbDi+S3DOOGOPVpjvHSHlc1UN
psmFrrkxJNigw/LOkcF/c1XzKo36i/I7Tr3niNnTnI0t+DkGF63stO3O41rUTmV3+Gmdz0RPHY9d
ovBzrbOF2/z4fXIqPHRylJ3Efd6pv2Ihyj2mTgzKYRcL8ZIQD/hCeczDrBbwCOfpPOUoVvlR8ZZn
+BKK0qWVUc26eYKw4BRydBfhhHngVGo6w2HNn2Gi2itxRF+E2ZcBU3W93D/QgSKFYnFkgSD0xjSj
oZr6SHirrund7hkmLMo1FzJDoem+SEu1aduD/BZr5IFws2as2NAti8XonaQj3eSJcJ9k6Pr+LRsX
9lctkarr+k7zMhjxS5ZB7Rqc85m/CuZQxWpc3rHgUchEW7XzOPes3e+H6VlKblVHquIa1kdAxuiH
AeQcQ1/typ7Q2pkd9TN2UPGIhjlUpSUwqI6GzOOjtpWtKCS0NDoMHMB2tFzUk8T+4AvJwji+lELG
ChRWAYU+UzXt6EXREaMZ1Jc6GZclINjDVV1S5c/JmhO5O6bVtfwlBpn3ZCcvFvDVKWCn3N0nEWvk
LdWFwwc1gB+0+FyqKyBAiSY7Moa6wiecwxrLwqnlQPOe8pD3Z9hKxsL0yCj1Q0iqwG3opebqH6Dr
uevTBHVi1PbTl08P7hkqmdXaUN0cfXUFcxNaFZad0ZSd6ddRy3reLuXP5Yt9rA4MdJjymb6M45pd
2hCVglXE//svm0/+OE0Zka8zivD4b/RDCUv0dtOkGgKeAsDuJ2F82IO8DLwfYxw8OevBLJ8R2wuH
EbJM5KtZebRrLLtFAZPvUF0QWf9NXQb4XX4WDqJegDksbxYEd51BZu6azInKEKvJGaXKsH3GtoVk
16t7474vVGKrz46+Y3zKCzOphpmXc7H7hq8Nibl0QCdqCwyD7o/bWj+4DernOZjxxy3IiikxgrDI
iZFbq31kEtr0Uzs3VwB2N1Zl4b4pt9yK/TQNHNlKUCAo7NTHvOTBuoRy0d7GdAQG7hfmCfz2EN+m
q7YSLqBy/RYMltYI8dp+L2W9yePe1Na+ZQgYl5fYMmt7Q365uuujYNZJiPPlEmHRdmBZ5W+fWsoU
yW7If4AKZ6QXAxqpmK1Zl4SRKwNZKrgVgIpKbUmRteG16iuIGph1VUa18di+gemv7xOMPSdV4M0n
Um/+JWnQxuhGuxcbrcqZTnfo0DPk5Hb603qpWz9bOnZCJR2lMQe2ok3gLVrKJ96NNzV6j1PrISdB
wkwR6/I4gsKPAAwVgQysoE2Qiic+djNU69rClv0zQyjj4aRO26rCcaDZndkg8n7fuE9kW7cHofyF
kN+loCWad50mGA4Yu2Po9V/ygxnjZ75PXsTDql7Sn6WqzXxYc6l3ZjORd4Z8uoEfq5WCBNKJHscL
QvqhDEqo22sLNkQ8Zynvaw83Xa5csvwND4+cJ8xSYR2hUCfA0t+sHyT2ZIsun0gY+ei45+5q3r7/
4tVQMk/lBIEoukWnewNzc7hyksVG+kPiODSpdqVJhCd9MlGkejGrCNyQgBvcqZ75wsBBB1yK2gqO
cVWA5t5kPDK7lEyXsHvrLAuKr4Oy1anJ66E8MFMLjfqcsNcGFjZmOIkfxDsGmit4scMNDzzb6yoO
XNeb/BhGaX1FkbHavs86Bjk7N1lG+wVQA/dhNg6k89+bNVV6iRyAbBhZWgxodJaRWrsbLJ7st7to
XFaWVtsDX//soNhe/U3ApV/5ZzG6MaQPrzSwwYyQ9Gt68vTP9oe0py0l/EBmnjTrFa7QFrH9FcCB
OuUz+JwqxsQh8zlzGEvql09Iw+u2MbP6XH9cVZi/pynB+PsxSen44zMmUF64VZzFx6P368yTra58
hjnvKWS6obFjCpOFeZh7eS33RLlYZj2fhBewsNw288K+1Hj4iNO+n4lUK5ELpwRWmbrn/1e0sfHF
QKRciCKtgc9plvvZPUcBfuYRWMCWmcv90BsKN7yu8AwNizzOuCd9u483zNSl7woTQrN7vknPIMnT
pls3Aj9uFQv53dtugRvnNthBKotFjgVzrKrNyLxXpjHRAPgKddz/Wikdxf2m9yGe9rhLovKpfMtg
1vVcf+Eq9BRJc9fDgBXJoJHCWB0CVOxm2Z91z1n4IosNXJTSwV6cP4gpzh7n9uUYUne/34MNUN0p
Kao+BbFkHMT8hR2OhDnYMSz9si7dCry9uEFSgXk6+bgMt/aJGdHLkhtMMEOdfcL2zw2RMjPny/XK
MEchlYbk1s0DVNRIILULX5lWmQSm1Y1OWMl9d+/FNx7GSbGoc7wAt4FepHGaB/jUmUFMGJ7/hQTu
cLUAau4VfZH+0W+fhw8JkoYeke2c1F84CKkut6L2DJhhg1BvGRZZEYSB1+d/8PUE8//Bm7olV5Ci
uVQCEzZrRYZsGmIBelelLZtHP6liX5aUMpReQ7zSLmF/O5tFbI4l5NVgkUEXA5zUXZ2WGCFC/5R5
H6m/4tZa4SuDocfArsEq6eC9TvfTN5qSMNkhkBOW+7d4wTocDNuqnneSocQH1s8Cds6IXlz9rZme
FpIFDSDlLyOjFDCbmPx1kRWvN2VnEasmudt5g4crqGAuUQ/F6Xn5Oiw7Ld+rozsR3yQvq/EkWoFp
aCdXFYFyDbzjYRElClJdhXZBAIzefEGdRF//vdfKglI6MTWdUE4liIRHXTB8iMbUG2uh0H4gGHS1
R6drMQ2TJJ082HZ8fla7Ezi/vQMF1OHIbt8bW0A7Z3l7a6wn6oy6Ndeh+3s100800d40MtkiPOYv
EzyU1wvE3qfUZ/ubcw+ATUmLyQ8mRoWZk9pl4lF6PAdjhbil9IbRvCMsKAk460D2m/QdPXJvM1lm
nVPsA36L2nfrsfRWFT5WbXguuFRA1Yw6/83xevmlEQl1NWKLDVI+snP6o8DxxPkVJFiZyL6qHpMf
zRThuXTAWf0Fb2wH8vBbHMJykwAVQe231lhuspCloTeA3V3djzqjCjzJ6jCdUuesPrr1SL7G7Hvo
E2drvYQCibuKjsuk5W40PpXVf4QjTQB+ChEKajK3Lk8s0qX1Hs7/LqAcKbF8JHtbhi/RdFbfJGfZ
I7JkWSACIxQzR6RKnc+i2dxoYGZ/BEZDOKOqPLQKfsNNMNMZz+Tc+YciKFRH6QncLt48Y/FAUjns
nMbM+7p4R49tE2IsRQYmOGsntG9hPOi2xIOYybcAwbPq/452iu4QDTTLSxuiFMJhY8hihgskGtHn
CqQY6roszG38pbZgTN7GjnBdSXdDxw/d5KwkSrbakinafX63f2M9e8lPzgzwe+9jbaXfsVKefr9C
l6OAHyDLzr9y4tjVKRjxFHnr6PoGkRQkP+Rcuf4I+xIgjl/ynhuDL7/5hwA7QIRFb1UqtnerAwbu
6Gi8ut0Yj+WddUGl/NUuDoSLAaL/a1V/oooIM4P4BbUEVZx90+KNpP1Qivds6Tw5a1sX08ZTGgkf
ZGWuFxkNWRe8pnxuiT4O/91tcLvlnSeoMnejeneEo0Y4p636fYpvU3D6hs66la6OgRg+me2PDwg/
Zv4I6pduUgnhgAA/C0hsYHq/9NodAhTSnwBunCGh6ckYWU/PQR9loY1oND18RADvpzVykMaklMi8
sBjQhvh6DOwiupAAf6KOmEmiy4sMPlZIrOwjMnBc1DpF8TaPBUl+H8XTUbmk/xXFDfHU42ntSnYU
WjXIU2nHaUAS36R1urAclCznanSHRuJDVRPUYhImsh7s+8/EtdVcxYe8rjdDDo1zg7MPIB+Hfj+8
7JUG9eD3S1xzEaZNN3+LMAIanw4LH7WV4T8bTBH8yvtBLjjSXKDLhXK1mSOqkxyPCL0iCT79oZog
GaoRIHObfF0CWmgNkPC+KfF13kYoVzsOj6AB7JM2p6a3aypBt0Y01tCMcVkx4laf0Og2laon60v4
y1yaoOauKW1Q5n51idYKZUOSqCQe0fWoGIxCmHZyDpUwsM7lVx8QcOJTx5IqxOIjhu2K7/ShIqJ0
K25XYd1hsD4AMt8Sufau2kiIK1S/QvZg/62efxCCJxXBYYVmSRA9LXy8LPJCw0OXScWq1ATJHv1D
99nVU9M3mAMYOMvudaskW25441+GtQlCVBexQi5W52fvbXSi+3iC+urvjUTg/N97CyqRhfcgOywd
bRi9C6QfQpLHaZg2o06swcI5V7+NSGtsCymggWjDnWS5RAPXiTdN3jottTTiMBYFoDjx8gFXlM+m
LLSenKfdPpLbVNqSDBP1itnYszZv6doQo3np1gF+S9lHchbR/yM7lY5z3oTOOdt+TeQFd1ZD0N5o
SZIRFTOYLWfU265RxBny5I35OcAE/1ziRlQf8gjorcJAqR8yBSuXeJ6KHlucL5Q+ZU+zAFh36+Ez
pBXbgAGMj8FaizgZWMIqZNVwn50ikG766bHf9Oy0V6CPSfDS5P3YpE4K/7f3Xq8cVYxkkqMw0EC/
AEu0hDm1b+9zvGO4tt/RdU3knPrAxlqf46Z9Y7nokeFiFhYaSyCtyhPn0O019DTNMIVjtlvLb8kP
TVrvyeA1gFoimGrt5udkFOUyam+DeZnyKY4S+rFZYyiFcAArBH0ifqzvTVVdIiVVKHhlcroLEA+Q
h/8mRYC6lk0spScrUO9+9n06slXybnbUiBX27BR6uxdW0Zp2oViAKc3HimlnbeqbTHPJ8mz6XaBa
FCVVoUU+ydntQ620mw3XtjMnGZ5onjzUlhvq6a91F+nCW4vhSnSMHAURPzGLeLb6s69x7NzyEEX0
mfZYHXsefAaPGGb7k83rkPzlhrOzkc2+rYhG6NZamlvIKzek/kmXYxh1yokzTfwk2JymefwGhFJh
FBUlDvlDc8fcEcO2PiWURKeM8jP12oPLk8TDoM4yZ+Mp4GrvDkSGg9KsfqxThQmcVlKlF+cxyUuj
vg65GwRYTAjnY/i2JJkEu7aaKEZUD0+OVvS60Xqu7gBjGEdXeRyEhDscO+Ica2zuZu+bT++Cax+z
hWRWuz6/9URfqK1ewU/Bz/78uBr0Gw8dXXG7ISl0dTdhifjyRWZq0StnDunRVe3Sk2YbgN6vmiiW
9r+JkvhmrC5/oyB5n9VDDuCp0Z1RlxTkuqcjhsWmCf6l/nWpA7AHtOOv+PDGLabPOb1La8VcJIDG
O3hXdKm7pP9A5uW//f2j1kqWR+ek5r1iP2yleacBsZMEZ921hALGyWWFTqVt8E3YJ41J67e18Fku
cxRrSR0uq6sYJ9M1gPLQiOVbp+Eya7lNGscNAVbO2P7KQOki5YgOPvNjRdqRTK4WwrYBzsAgglY7
xLM01gUOs2F+DLyKIw1/FKptwsHGi9BcysLc/9pzcB3INDs/51zp2XugLQJmBVUml8hN2z8LXb4F
CiL2IV+aiHEIfkW2s1F5IQyG9CWAeNmHluy1tQLhx7TE30ZVhCO5jGnlhonz2jc4hbsTqCfRmiEk
CBe1UDa/SohXyP4kkn7u9erSqR0O0rGQzojz74YGSO4oL3IdHNFl5shWOLyI8HzcEfv085/2rlr/
JBJ7spBblvKVxbu5GwEkty8J9408eD3WG5FZakllCSYbsZi9bI+CEyUq0uTQ8lWVZmya8fxGPB61
T4pMq+EhiSv7b/x5tUMPOXQnod9bvBn9e80sLRhhTVS+NfU+byG00TiQ65Pi1Xofy2Nrqk4+CAaq
YNcshdAyFotT8DSXwbUcS4ZUmfZgICTlnTjEyXfji/c1HpIwjP+nxi69tvyPHmei3D0cwYKXkMnA
gSCVBiJiSfLuB/avQLNaalpQAtjgLMrnruAaVVz8oW3gjtBWzKEPrqVMan6u4+QEi86kGTNlgYXY
YwBnYyDPR/jv/74TZoSKr0AVtLSn2FJ5dJFpZQ/6Npah+GYUgLAMNvq9RlknYxppsZa6j8NHm7VF
uJvOAUGVYB2+CLceqwTloH9czP6FIvLQuuI3L8e2VeIKajUHSVEDzFDg16nZmsEQM9xsg8KtoZRF
iCpQK2VUoOAFWai221B6sBbvOJKZ9hibZT8Vfq0XgTb5oPABeVTZj5w8YBrF0h7ZmvmmHarpZxIX
KHctA5cgTUdMZanT0NsA0NaFjn88OkJrJ+b7FWSIAMcXGkR2xCrMi0UbQsrWL5CHf4eZ8TaDOyex
nvZh7IZaCDZ6/FvK0sbb72eZ9ou/HJi+Q2ENT1QI9VqHp0C080NHC/VwFuhlzbAbiRR7FadVLwC1
vKczix7+r4qa7pavqMHSXZjF02MbCVV/708GMXpUmYSaiqSp/ZZG0PrrOOEealXN8jqY6U2sW9uZ
qA7BjEbHZPwnaPXac6HyYLq3mC8iOjkGD620EswdcHSbkt+B04hHNtkIvn6517hKXRjOsTQJj0lR
Oa2490kemq/cGjXlmSQCslCPhYQuMIlg8NUQGCWQRLLemeQ6tfr9iFdBa+LIY0LXTngJFsBt95Wg
So75czy9kzEPGDsEH0haMqDZxDq9iCpIXzO8gDQTNXaA5BDI+5sU9Ni8sCmmu3WJSkUwED/QFgd5
p4SlYYA7SSRvCURXoNwcJ9WmSZo4tgOATIMlQynXrLCMRj8qoZQkgSID48Zpx5lOBV6pZLtXmX89
aQIsI9Mg7Q881Jk3cFWEeoinRJnwmtc67Ova8TOHbK1aSnAGdEYzJlyq0/cFdSaSIFxU+PTsrllJ
O/pFJDfke84FfnNfNu5XmCYD0Ggq3IqJ9AQHLUg58JCkCLPPuMvmx69PltyJhmq7OewpqNPeannT
IB35kWMfEEo8wpBZnYOs1WIUEWqIEXyT51bKON4gIueaZWRNKjONfiSrzmiaGe51LsjkXmUtf3zJ
sizgfmuAWRIrwAimrctYI59OGhJZNZcjyjW18Fwz5CEPcg2YLtVBAoNrhbUc/5yYVz/EjmBnOVgV
663sq9BvV5pd3VnKmeSYhtTfr2UtLmXpygXC0nuxrMABjuvcQNSRKOSGysSAZW+05YDlzWp7pp/R
bICAwfypsg6Cj0oIbyBX8nbTakZfUWbXkYPjOeU5FzCxz2joJfgazqz2IbX2HW864dDLRghU5iBx
0Eayv0zQ3FEVJ5WGfebBq3GOcbcdnYtRNd4gTCKyPqvcoHxMOXnSCUygLtKQRzqscbX3qjSENYg+
bjukpDmKJWaU9UWYaFjESyI6zH/zmpeqsPlacgm3wkeRZoEw1po6BadVh+FqFnp+G49z1bhfoN0q
o6R4qyuiR/T07hUT5V8SV1GdYznCV8wMkl6d04j4s5jY6oVdbzljwHWzpuH8SSUNL0BralD0IkyK
kd6knIcH0lQLpHtjI0IMkR0JmEq/Lrv5AqT0mU11k4amn1UHfin9qhVnlTFrWqaR+YplEEzAMiyi
RMRtJUdRB3IMqFnARla+kFYKjRYxwimpc6i5WLOpjOKb3XVfcyphcgd54kwqTzOiqRvr+/MoXkyb
VdRqLc95GulNMjteW3f7hyiRCuOW8AJVkPbMjOUJJCTpJ7OHzbS+xwBOd3TF/PMsPMk/WXQskvKz
atI0PvJG/5+ierYxzGGLGAiR6kH2eS+eVnXhuP6NspDlwYpS8jL/rc8TcqbgMwMFe5ZA448oBxM+
RvRXLNhHIIKAHXIHxy/6V6wA7h8scnpUDWl08jE5QJPoI8QX3X8x0tMHKy88/TeqZynCeUGDqpa8
tShA/vVH9ktzRHL4MkMPFAEjRPSB7+grfU/TqsY/k1Ej7UOfJwQ6GrBz1miPJGGbDFhjB8RVTaYF
DAkgZaliBnj7ZneWcvSwVKjrgnKR216tFGJTRAuwZgtKA6o6g1x90jcK2EoBPphzmWQ9UzP66hdA
Z/qx2R9tc8Ppz1CyCDbOWlLmWfoYIK7QYcFT5/L9lb+fJlHoZuPZilh1TKRsXhFnT9lS64gCklLR
6U5owjOXJCvpNDcHq7S8Rvks1e/yG6g5lcbzyMwrQ5sAyXOoJOID0gBw7UrwPF1vuXcfICXchekR
EIQFVs6kc6sv0yKcxjIyh20FCnWRDDRWEO3K7EC8i09ZI7zgBqOpfLeEVB3X+hjviz/UhwkjSZfE
i8EDPLHCVATEWQSf3EVlEd2lHEBucLoGu2dygb25VtWUqUG2xVbbLjRIlLjlbPuyqRV/rwzWbhjc
8LZhPhE60uS4YVOBD/R0L7aHFGqNSAfTBG+vIjp3IyYfr5qMdwgOOr4T0eqbMrkAdyXYg0L2tJ2O
N/AQrQIQfXhefg8dIFieKswI9JFjGuKfPmlAkxQWolwx9QQgV1SCpHBQnr+5skgokoR/DhGxbLOs
Q3uvAbAPWvtgSHAQYuzvPJ570IZvmoz8KQ1WbUgWHI6lwpgQqH4PGNqplFt58/Sg+roNBwseBCsm
wOzalA41B/rvlMyIAQmm/JqXmr6j0yPZKDNJTXMz1Rbi9oexzN0DXtq1bZw18LUzfR/uBOkjPp0R
qiFKapChWl6Q/jK+Hrn0xlh6jaFbKe5FGMQ2WeYcOh8IdTQphjU2895hcDT790fN7PUqzHTko3fA
oy+nLEiC8vJEnEzOsVqWT7RpX73nW0OqeaWghNuaQEFGwv66jgXik7Q1XqezHS5jHdaJQbXx6Wpm
+NKfFnueO+OyUqjfS4NRC1ky8rW+Jaffa/OwXVjOv8YCL6MLRztt7oXMyL6AY0wsOlfz9fm6rAt3
348IXrhpghQgMcjUiUzW3DkyGIj+Ar+XoeTLG55Gf26U033ZoFJX+iAUzavpwqKH6t+UtERoJjms
2l1S0Xy+5Qh6JXW9jByON5b2crwCiPazL1dd1liBayz8Wwh05cvYEJ92x70rtOcm/em3Y8dO3QnL
F5YFLDChKPa9Kn2HVQ9+M9gu2KukwC3NBWYJ2lAjuAb7maeB5XmEqYzmCOR9/nOruW0vHELFMFBr
Do5l7PJFX8TbYyTlAGu4nuRgKtBREAMkV2yPEcUgZ/XI+WXXtojkV1OzsNdOARaw5VTqQdvmQ9Oc
tRPJjUq6iO+xAkX2YE/pTncODBL5fPrCqyWhUPgh+8sD42O5WlZQVh8MGmGFtOYdYxrcLev8m/A5
FkW7656uS7UwSVsVaD9XdH+GpuIJKlAxJAcnNyzwn7wU0wMlUvH81uMbsKNXLVjitOSPDEt49wHt
/bOWfZjxZcvqPH8i63CUNhCNmkeyTQgjvrkOTPpHCKyk3enIZO40AuokSykbz9WyHgWBAtNQ67tO
2j+1H3a+7aVdKI/026isUVtp2V9gC/dQD73stP2qTQD200rNxz1+prEj/jaRZRxinwt1jA4PU0IQ
gSqkuywHos6JGWlNs6XkRJ6LbwAVGC8QqRNl4OVM4kZGS8Ls1GyuavmUUH+DrDMKZUxFZVTHdfrL
jQPUuSI5QhbY3kCFOaDmdbbha3DOHhkXP+qj3p7xre5d6zrmz09pZts6FIwtocQ4+cf6p8yanzIx
CGMCTgLNlYK0ajGqARgbmYHan4Cj9QFlZGtO6Snu4xHZAepAC/RKIDAHqZmLKeQH067YiJgleR/c
DZ98x7YRUxTTIdm2szfs+OmifSY9Z2BYjM6cb1b+Lp46NduUTL2BYwSJj1umdUrZPFw9raqVEpVt
CzM+WJgFhsqUO0notQQ9li5OFWSnPE0P8yChIHyJqwQw0g/cZpq7aXD9HCQP370pXHQBI2DtdFXS
dYXXy5ElmBf+7+Wmhf4n8pySX/h/Aaf+eSkgj2N5NbSVOOAQjtBYkD/BxrrNQRyrPQS9eEiJjgRV
+y3SFEUaDFN60XWUPL4PU6GpNg7pufRqlwQzP9UGl6XKwCmh7UOUrbuSplJJ1srTCk8b5/yNY6So
1iYpd+gE6Ecf6TU7MZ9lO3g26dadJ11LZrx8h85UPoXc9hh88jVQpmy3sohwWL/sGGG7bViGL6/I
T3Zcp8Q9yHAveyIfZbyOB1qkPLC2xauFofNIB/lqq9Bx/eeObd/mA0eN5Xea6ribPnqfgizqt+mW
1OictD8uTozAZbuutsz9uAXHLAC2mBuZidrSAbz5ZAB7XOwmHg4S+NRzCE+aZOhnclAZPXCrGNUX
7RhepLS4h0sLc9+kzXRSILDqZcXJ33LlJx/tCetolWrXlAvx197yJVRe+0RY/HqCZ5+JdA+2Q9cy
TKxc5AM9Vgy9LD4gfSwzAbfhM8XzVBlV6qttrUmgmWHPmVqIYbpHoTAYDtVRYzKIVESiP9tlFGtR
i3YuTBgmW3ah80LfLhLlDVwNGPMTKJofXM5nHIumZypbvxOjI8mc3tvisUjh4EwQ2jFxKRH9McwU
vW7rhb+Dz/oN9w9PMIByD0UW7ihi4aFN/YWbSmufVoq89laKRv9qsznQewayYNaNDqTnKx3X2m0a
9fPPjOytXnIEN9gA+A0gcqw8fEAmgwQ0QF+G/ZXppwiaU5CSdh8JB+4fTRVZ283RRTD+1Rqqun/W
n1nL7NgrwLDN8sPvSi5pEtb0u51wvuSYqLlgsqlWNIXySUN1aAWNXmwlO/rdOQg/j6v3mJ7zEuHm
dWPlJAhYzDMVt9TUxik9BUiVzPCOdHlaY1a8AkrbC8cYeXYOD3B+5tFp8HRJqSfkrfZrX8OziEXy
NteuelJDaeyyEZqFR92GRXAqbmlYqNlZTBeGHU6Km1E5kxY7looifdZ70LgUrATHJR8Z2BcjDI3E
ikvZovqTpuoW8LzEJYV6NJ/futot0KvyA9kKOjegvN//CZeLa8IAaOW6yakKvgVBPTuuMbO/XYzZ
Mtn1+tkwVg4P1tyfqZ43y2XPNpiEEaadU31enSo21ID5VWqBxS2E1SzcSrb30N6rSwH948z+v0rH
PAPc4bl4AhBL/Smggp8aHcatgGV+/SlY/YPyUvhyqW7LFyADUz2ayLGyFGdbTXiT2w07d8h6Ok4Z
+BWyEw6cezE6SpwWK77Td0XpJ2K1ZvFtyxuOOS7ik7iio6ts+QIaw3yM69zS59KaN69ChAR3L3Zo
2PXQyAk0MOtDKmXw+yclOeosKeYwRbGHsf+PPTVlYDzaiTLGAkZJ3raoRnZ1KloF5+lEObPt0XOF
mlH5+yvm8Be/0plV52pzu3v6TklC3P/3Pki/EFIGK1T0jEsbqwWw68bb05gSvIXXNMjX/33pQ6qm
E2RZ+rjkcWeNXUSKW71TOc1OQVxq886r0ULWW8FyC1zVaALQVZQITr5SX2hQQy0ff5G+OZjseDdS
JP/sh9R8GxkPAmgiKZCi8pJ7FKemoZmU5iQDr9eS7stUo/zrKIYTzefH6yeNaCgecG28tLpPA34I
7Bvhc4pCX8Re6NnsdMurdh6/ea4qYskKhDqWBUFbRQl3S5pCrVjun11uI6xdg1LwZEdkFOCWUrye
9hoHdI+wznKi3KfbRIBA+hg3jKTaS80zOSIQDLHd1tnaAx9GwcqWtNW0clXqu2QV76CasTp0yRmP
hWceP5MUyXAAvhhnRJw4iR9pZkztaCnj9LgUPyMW9JQAx8OgWN5dOhV9jUjFULYkki/9tkx6NPxM
DjXIQW7kES18DglxzHl0Y/esErh1n5GS36iI5hu2SsZeUThTLJoaIhGKoX6b7v5EIvNnKIQh8Wfw
Ji80D74UVSHGlsisENfZ+51auRIKOYhxLiiQpxW43FqQf0qpz2T9NOm7oouC9uQ3j4AfCPYl2X9j
ZDhu08Isiha93tscbmTTDLY6PtGdE0tnLJLwCc2cpaupsU9UMGT66EBFAfyyQiFbIC+AsH0yCGCa
GhKvjXM4XKAwX5f5njNFLibLYvdTnhkN9HGtzMqOQ8c1TMLa0qtPbVMKk41WHAA2z4eIEUSGhi2T
U25ZIl64aWjDEVo12eNc7ljSaG3N268QtRm7/ZqspyDNvU8U5ZLiWnQwn17q5/O8AIT/YO48IWJD
t2f+4NlmGKp6ExKr1CpjZMDiYbdikg7acDZIFbbHFRAWr1Jv8nTaJ4jpr3ozmj/FTb1QB+bGl2Tt
CXmWo+6cHYH256+ce82IlLCTynUpEZIxFf0mSijJF8XJzjyJfQHDUF+fWseIU5mgoXrgISPde7PT
EzFBkwIrDz9z3twtShVqaQjLk6z73ye8uwFNnICoHxYFXRxpSMxql1RgzFWnj3qU1H0yQ0pZu0Tk
hWvQuCi6zigTZ2DT3OstywGYOFB6xLDs5diJh54ol6EDLrwz6+htpH6Slq00+JSut6CCEQCshYs3
Zx/gNSt4m3+h2krtv/e8HCk1zTl3RbiZEApF8JBhxmx5OTbS/6l8I8gfi5U/oVVpoa8GDkl2B1ww
Uz6UJEy1xy2mEMdJh3s2gAY/qHaSIERRI6z5Xxg6C4soeOS1Hxv7FZEj94RIJnA5a6f0eYGpJUSb
n5uXCA5C00AQ1AmnHtbtJulrAAbuOBWyVA+UnKhUyC4uTNhA6kHJaNYDz+7EzX9/BPQnXutDuBxt
BOK+bH1Aac2X7twZb3MqN1nyPZYRxwe7Sob9xD3yudcxxFmYshtQTmTZaLxNku0o6OYVE5U7zq50
5PaI/VpwpiESAw7riZYua2PDT8g4fVp9JPMsNcDRYv3qKzVerI3fgzqq0x1c40IqepZLDFEHu6EB
gB8L2q06BewSNLg32x4U941WvL4jhI4EK6n1sXF3Ru0ngwYgb+28iAHVnwQL143IMXtkGjmSXBM2
CvNTGSNfMYp7AUPFrtUiK/p1pGCXSgRBRdge+UjfV80yB2gYPd+SvJVP8RgygXI6WYY7XsCNC4iB
tG+sW8JXsU4ugCrnaj1ZdXRXanyc99ekAQv4cn5iQBUp0GlTshsiEH2zeR/VIWP4cuipIVEs1sEt
shRWWebLcXTSG2lVBO/TmflehdO+I0p8B/hH81JkOYe9JKei+aJrgdRmqIZaJOaUF+bP0zxYPh56
Dl+1vPSUrId805vS/SimMzAlPJcm7zUIC8gTR01H0wRn0FcRZVUHdMWOFrmtw9wUC4sZsWELTyp+
6v+SpuTXoiileBgToiusOVky6x3plSwcLpcMkRfNVwbjkiso2mat8bTWZAvOGY5jldg7s0RC8qIr
pdNZ/E3ir5fSiUivGuCO8DdVu2v4Frgc/eXk1MwXHJnw+NIrw00nQJ7nJNvqvJ1UMDVUtEnW5dbY
mrBCk7X6+QfikkcDMkaYORobYTO0g/dAgxASNj0oLSbIed3Mt+IkhrAa4ciuhjQfMSDTi7BSBBTD
VCEP/2NhmO2jIbB54iNvnaUXMT6EZTxh2EfBnJ/yy4AYVijlAsLPc+StvwAgCDIyWRqZ4sosGGpH
QyYMWX+PcBjv/1IC9YBle7K3TFX3L+KBhWc+QGhnwsiOowFqPPFI+o5pGz7xLQOyYwuJlqVeLKhK
/cG04gmnhzU4vSj/sn0CFpRN+dCfq8M2bbJsQKPYiCmuvDalTrH0Amuixn0iOoM96cACHeOFCCKP
J8P9XdjWUdc/tEk9MnEqVw5fazKogAkJVZTki5kgWVfSzUiTOFQDpagt5kpsaX/o3pjq4trzowLo
2tjx2kizaVg8khVG4DURGRMYkx5lBBvTGk4tOWv9cZ+zJN7osrTOCANqslPG8kUk17VpMEo+0kX1
I1Epe/4HgzuvR/Cz8IRNNTJdlPFt47A2F2macjNd9Dc/9rRX/tMDLYSyGEEiHTBTb7DYNUFqHMoY
Dr+HOWmW0fN08ObmN9YvfRz2dEfhdDYH2Ma3gfPzmgigqt6Rhbl5ZyQGqEHSacnuMmzRgZ87Q6wc
IPxrdrVBzkehYOsTtmy5FAUmyI1/rryBIoGHFTMqA3wZXAkfJhOBEV2biJBWQN28C19p/6USFw6H
StLJqSEov04FpEOHxXUyV7DeMbgn2N/B3oLeIH3bLFO6cIw10jKiz5nyt0eqSzNNmvXFCfVRxNhH
ajp3IH05tmlGHQxCOvoXIo1F6SdDvJ8U33bDlBCUl0SwfVoW4Ta2P2HvrbkCTdatEBNq/6vqhAWM
xLfEEzJt+HM5oee3rpMi8r5p4nJ9nGNeBJcJNtn4RtAq0gqzClnpK9dxlLH9azrBWmx/gWERrbKl
IWl6WS9LG+sozK4VhYL2OounNmjg4SlD2x5kIixJNnqzydXpgQKRxyQjHktCxJQddFP1MziI6aHD
Urt7HyELJVsBTqXgoZ83aO7dGtb9f0itgDs3bPSldFwAMtK3peLVyiwrT5QlJEOsS0tB6JPE4BTq
YKPHl/uJnRNjUEZj+jcDMN37QovxkjXCilPg7Wylbfdaz9nMLW89MACAyZiohFG0ZH/D8qLXTkHO
uUSBa8aMVKbigdAFpdGn+zrV9kMPPojRFNC3OxtOR9+kbhwfBgwZAhzHO9EBhQUF8DDjHAQ1xLc6
VPNgaw/xPIt3zZVvdetUkBHXo2MtPOxALRJk5s4wJNpf4lDI+H+IUBMK9skZno7+/pIFFRCy/f1j
D0xLx8/sG1s7hHAw9N6Uec9l0rDHaLGXb+PPlXuQN4EGbB/WHbNwZ4vjGvPvO2Baf6WD7RvuomxG
c/z/GPhmrondYck0BQ3fqHAtvCo1VNnZfqrYyXRu0Xu/MqkPMqcV9np7giZkpfO1ZegjmapyXNtN
x/ay6ZZIpMRu1g1oClnlcV/y8hqH3gzXMdl3FDNfE8cumLuzsvI9Mg+YH48qMq65j+3GO/MpkmJJ
ONUvJWHl4V//EmqO/pn7z2TcwbpcnDrq5QyXyh1iyUw4mon82uQdHdtXU5dextMx+mDhQ0D5yzK6
1BaDlE6koHeEcNSKhwme0SzSs7PbJr3+YklNH4CX1B6yk5Bz58Iyk9JhqD5xGKnKlt5AK9ALMywt
/2dMRcnrgKywNv6CxujnZJI3Uzmz/i24YdCFkVy5Xjheva9+YCGvxkBS/EVYQcYDRl6NgBf7fMZE
AbM9GMUL3o6IfyXAoX8i4mNwlLAaXZPrW1Moda/qu7UYlqOep0KVGZhSo7ezO5xZas9vsBV40qUa
JKHFqp+hcHBp30YvGo2UpW+J44DYEXDqVLFxZ75YJJEJj/RqnaNyzBFRk7RdVaoRvY+bv9G7Dv+u
WfAn+jwtwdHd/2vvL6A93LUAZDB6zIOQ7Pjki+Eu+7dm25gCvp6E38nCGzKMP3RvBssyShJkp6GQ
THebk6DB4djViZcbaVxinSOLdh6rdahQJ40+zG/E7BIdi2ZT9jokKb1GTxDrzOvUVh73Wnr/Oj6C
eixiGkS5Rw9eFBPaWlk+ZA5kY5hfIWhB2o3OF73+0n8BueUj9uZH4VWehKc46EvLXD80V8swkGsM
/Zin+5vQB+bH0LctZtz1vnS03EUhtj2nszQACqHWbNxJEfHQUQttfNFax/TOFLvvj1H1g6YHgJzz
Agfml4IRm3vKtmmyiY5vUMGDINEqiMOi/xyHLr/wsZPZbjjsMJLn/H1gLMgVquJIEI4vEJsmxpHW
BzV25Cr2VioFnN7UEn3S4X7UO3Ws7R6gzvXa3iLiv4afj8+4DKUPnPOrg1MJiGWCmUkdPhMO3ReU
mu7GMK4wLoTD6gBKoOJF/Gh4HMOLDYZiOX+Y5R2Cd3ptKCh90NSprJB+ScNpKupGQ/C6iRQ3OLBo
XoN7FUg0ujv+P/MOCYx+wCWnYqD286T73rpwx6jwtDgUGY5dgT8zjWyskivDzSusF3Zd0gpVEMmp
NEdNRdFPqh4wRwbmJVH6q/loiNdzBtDvyvlB927rjXv8wbnOiMHbNb5RxwCEe8+AT+APwpP41xZw
xQMKU1EsvvV+zJfo2oOizhye1+UayW27v0A2oZmkg9u+frRAy7id8XmcUHOWXtb60qSSrSWe82SM
9rTmlqqHx4Xrc28SCA19LLm9gND/UKjNtpmyMmO2RUiluq+WqOU8EsZHCgwdXOF2UVh8WBiAGmRn
HzSy4/MaVrGjk6FWBMFRyL+s/Z3vLfmkZXY85Jo+dT5LiheA59fdDRf1iE32jsfYqLn6q6PVAast
Y4BUNYvTjH9BfwYwPcuPvioBDMkQJYoRh0HASACLqsrTXB0ZaqT7N2kHhenLYtB/rBGVgwmq7m/s
BYstjh9nSr4gkAbhNo3A6vWzqpi8Wr3RIgWFZRiZlH92iXTnPD/JQftrypnS1aEQDeKLivJuIzMV
ql6AISLgK0eUAHiMeyXVl8phaDvTilHCAKtvyqdySQRBBQ9xwOItfwrKVqwlNLJ9F4CbQaYRk1Yw
YZTeS7ASrdssvDm+1aGbx+SCen4m5oEQ7o2MdSyx3viDVDq7/gqE61PxJbQ9O0tfHLFR+KFnYL5d
OAoimxLW1bWs3S+zBct7LJbinpX3KkXhOcEzY6CrDG2PxnnyO+NEHCdUueXSRJaeCaf1aihbZAQM
ToAS0ZPLKxoO4BdrqY2lUiPMCvMF37L6YrQuTQAXr0vLTE5y9tA1PmRn5A797yKy4fUwQ/aJjiS1
APIq+FWIi5pkRDlG/UoeCWmyx3kFyA1r/tUgas5miDCIkACcT5BmR6BdLffjMjHFU8SY3lTsSfny
9FGT+BTugVSMLVioYMewJv7JeFRO5nEMlVoOCZS1ZYe5M/G+KgMSD4a3tA5toG+zYx4FS9MrYWJY
4s0IEczJhA0usEFOiLRHWp2i5m03LD/MCYcPzFfYEW0xLlX77wY5QRtoOoYo03mV+uIEzv2cuI+l
v3BErv6TsRSD5Tl8Y1a+ZThMYbHjdBb8M7C4luQBpeQ4AVQ25lAqk8hspr5ZW7rZNLhYOwmDduQS
USeYbDKY7vDXQSfOHV1TAx7GJsuJSLTcfd1JS4VSNB0MjoI8weZLNN7r0+umJYTI/CuY5hgO3ygP
JOJg+Hi5FO+T2pyCcrCxHgOu5pJXS2dl5nOg62VQRBaalVQs8sU+WaaqBfSxPo0ZpfSJOdnynOiD
bYLIYi2bcvbeL6Vy0+1hy2YM7qZNuvUPuyK1IOMOV+oWqgr7ad5MnS8FeE5n1Bw/sn2hvPrPbqln
mASwC/wIzVgb/jGKKCwEyJ3edzEpc4/yeYvVGsrj27w2B2JvEI+I8jOyh4HsVWTrWDUFQy3VUXkJ
vOmic3xZcGxBz7QOq3dn2/KzpM/OL8Stl3j8aX9QjXdQ9Dn8eez9nqgEwF3TFQszdZYCi0J61NNm
GlTfngA/5teJID8pQPuMsIcgJFdqVf7HpJHFx1dA0Wg1L5zMbpQqzgIvEBQ1I6OMkYqBSVd6ZMKD
xX36mIAp+prAzknA6fc/pQsSHvmps26k6Fc5JWcNqTNC3TtHF2yOXSxodiqd8/Ao+fuFFjJNt/N1
6S8PyslB+wxycOSDhf7iF3VwxR2ZNkj6bRJfj+Bpp58mDUWJ56auHHIq4WsT9OnuY+q3Qq/1+LTH
xPPU4OcVNCoFUcrfHXZZUne5P+kXyizzCaE0Kz+3ULiPKwN/WAHLFcQC+khMf5Gm7ctzPnR2h09F
+uu0Pl302N5QDuKlYilJVHkaM14aijCYAU6HGuMORbAlCcdEWWmNVjzEMYXN1tpuWIjdBX+/ZZiy
PzoXDAeE50fgo+hAakqJCloWIqW8pAcv7zZScRee7d1nGw8NtUfC8BqSnJQUC31rjPcOW6hxgRTJ
+AstlLejnSWhrDNfxN8KFCv3DNIZUij+ZjvjSac0jZlBBRqy5KEPTqdVKVYfj33glcx2qu7RvQmC
vDc2pk1Ifgm4Xp3YEfSymoMvtKDc8HKoDXB/7lIkraUVV9Uk6KNC32a+Q/VHnQu24kAhs0t4YRaC
MhBRTwUjJNhBmwTmMCECeTi5NPkXI8r2Wkuavrt4O7NNjD8t59SK3YvT0ZKdVcTvhxg2e+Fu8SnO
7wAUbi5CtAQNID2CB1Z3Bw/9obE/mMC/S3C0rL0VzOC8iWKAZP/REucYXn6WpKLbJaxA8H2HB4Sz
TCd0WJVAO3YwlPbvfsCzzFqp6gtkFIpHfAW+w1wKgq5yGrkP2xPaN9vL1XzFotncSXT929xbStym
NKivHJ8ZbkGKm65iOCtNXsbJCcfKbcmEg6Z86zr4TGzctYmuqeO5RxC3cODHaht9CVAVe+HGqQdU
8sjUsoazvHimv2x8/dz+oJPNRAXPbGWZSSSoFn0oQZn27xsR7cQuG9QVPaiSDWbp8Bb8c3MHi1s0
mrCOqPwUTQGf+K3t8GXPsoYXkkZdOKfK9hI6NV3q2JB8Lv1QE6h0FoYRs1bg8PXST0HJ4U51DpJD
NObkD/OHaGCPekeqj6IBNSNuB+y8BMNWXwhkCRSJBaBtJAEcKuXbWq5xDwAwSrr2omLv1Emq9DKn
U1dEbnH1iFL0SAYkO5IhQl6xU0ulGtmEKLyOWUpwVEuG8omGMUyfW3aNT3TtJorSYR+9rFzFivIJ
TC8/y0n0kwT3w9uKMkFcBflEtpCe1psLpxRSlIW2OjH+dbUilnv9UL2yp0CxGn+yBOS9HW9r2Gmc
DYH7UcP4W+w329+06kQoXFUhxqC00Hx658eh3kIIRzsTlm9WfSq6P0eJu39dNuZ46LKpNw53ec9F
VKqTWpPzsNEn9HK6yGpFixDxc4EbzIZuooeciBlM7EBgpzHc7OJkG2lK6vSDyjIUySkeIyV/UyAs
geypNoudPqgkxIv+Z5Gz2Tg/pYvEk2VyeXWwnpXVqy12TrEIHmkhoX8J+S0rAmK3aSHGBOAFfuT7
ibnNjUphExXrsMXHEBvof0H2MuFXx1NNVLMP8xebm12rGH+pQHEWLlohOZSorogyJQrOfgzlp4tg
xgRISveGz+cca1hdzX9oTURYaGwVaplAnygTQ99C3fouLc/KUZCFLh1DKqYQfO9fL7eWEvFZpkyc
4bNV0jteCTeDQhdwY80Zw9saMQQvDVO4dTEXAqIOST0tx4aauREb2BzRxCevRtFyF9CPgDZ4j33T
h8lYHefs8zTyaYscaX6yyTT5icLoUCl3TMzjD6X3xbD5VptwRqMU2I2ckAJeMgF4WdPxlLUOlEhw
BpGoFvyyn2MLR4sBfaybQNMPeLHmLV7jTANVKSt9wT2oSvIJJqmf3oe40YIQz+91sBkHCrcnm6za
B7fynMx6fr+B1YV/7xmrJt6RsKy0oCIVipQZ+rYA7H5lKX7pd8ykW0z5ZlgB6kireA4uFf9egGO5
mloK7UQi9NArlTz6+LScGnPeiaH8WngLDti4dubk4pXEU6s5gubb1tXwphXvVYFccbVf8exdJd0k
kOgEKeqroSJAd8+rkwbhLm2UXzGHHY1PyaZJqkEF3SCvZiqTjQExoSqbvgUvGBfJuy2I8xh4mP2N
BT+RQYXdxxneUzda6aVmH5cE2bcOfntEd9VnvVMIBoCTNI+FdDYFUFxzDdHctpTA1/2+QZOxNCeV
pKMIpI0+BZyOy/AKcWUTR32aNaThV5ZHvSHbsCXoCvB0K7iQ5nz0mlUJsc4Ha/fCIOP/B9G9V2GY
hQbZJrX5eVuc8uC+uhN/Nh9X6vPnaQA9/ysyc6GNaHYOl7rzad4i1ZpJQv1DaswdwL+TXIK78gNS
HZYqeriYMMMKX1wA6lixwWX1EblZNGrsLiMk2Xc+MKGetdJP87ZsZul9rOjv2VFZP7aKI0bHTllq
v45K8VN9toh8u23LkPAZZopv+XHMP7fzoKjH2fQV4NwCXt8a9tqEQQxRA1hRk/wW8qpB3mfvn89u
0/b6ZIstlQBWgoAtficrJeoXw6jGkjkhNR8nW6X6IZAjzGaLyTIev+rmK7b8HbOvHDO3qLnj7I8h
ct6qskcpsufecV7hjc0xKjBe4kau3Qxj7f9dULHbUS4D2kTt6lwcHQ/gKtVeZhez3VQE/lyS0R7p
cUh779BZK5umPbr610I6kMV0byOMz5QTJSxyBt+3xFTivXWHewsuOgWoqaTCescudwbpnzaP8/BK
WAD1YNOb8TB22zJEX19Se7bPe7RZpNuPasG4hoWSQAOhNL4+ZLfTH658skRGmPvhtvJFNkcNLr0D
Gp3Y/J7JyEcfqouzC4jN81ASJq+SvHGVVKkWelp7ZnhWgRMVjtcWTpEV4iBJutAxVlxpJOMx7Ixs
hygvxAG2bAUH6H7vI6Ib3Zle0jpTmGSWMrOVbz4xXadSq9SV0iULxgcu/TkrDh/mw2sVZR4GBYVi
9ZZBUTuLuqr0Q0/swidGqmuxmLhTw2QnHxCuYow04OUbfnQmzNFr0+j+51u7l+00yjxGcsuKVF+0
EMGUKccIkN6+8OORlnqQXSTZ2vLVgn4X+nc0ClvJexffy8N6ErB7SHzOyfV4kljmAzXwd92hXYnU
8NWgwICJkpk+ZZ5gL/FxOq3NRlboiF4+rKRT7QBzfLe4zYgrQqOWc0Xu39m4jx6T9I6xcjP0T3yo
pQl/qWvbjzfNtxQmaZy5rgsA0TKYpSD0H6M9rYTw7iKt9mv06l/9rlxZAV7ypZn59xYMzbCKT+dI
JdYonOJwctFVkKmUcs8tyPZwnAXASI4NpRm0AooQwi0Ix7vDfSNOB5jJW01hVt7iwgUpZavcLlrw
N2AiMEG5s9zlYhjzwCUpPHzr0aODTD4/fzToynG4bN/SIYQGqcen4VKSJGMk33cjTCSRQcJrllbP
07lCFfRn+tw9UHn3nEpRt7GtwPS9sHFC4wP/XreIhcWMfkBjgfRcxqx8aab1OeR3rsZTrRibBHUk
XCHnf5x/x9aE+GMyP+PfoAiJeaap8tgT8ezhjZGtlWYWFTSqITrz7U4EwdzLLFk5aUOzR42mNgKw
fSCsSpHK4LYO4WxWDsxjA27RcHhQ6WKgOEGBhJRvVonn6zDa4/WnF019BZRjcLVSG32JcsSpMrAl
I9qrN9AWWCvytwwyaShDK57hIhuBQpTLnBgTAKUTkMw6Q8mH8mT1+q8PkzhF8FAO9D5e+u5cMLTr
AhqT1Hc7uSgQixBaLjbtF7g21QorpvEo64lsLLUyJSk4fj9H8wDwXRBXoXyqkGPpswgDQMT9QVUc
nWm7EYjR2aagFpqirlw0kLiLrAWw1P7oTTp9+uo6HQEI5+9TqcIlVe72DkcaYXudq4wf/35nmy3h
D+3UmzwrBSQVT7jU+hPk1uPGvpks344nvE+IId9sACYB45aN/B6BCH+dow5G7skTInLUDMNFPYrr
rDCPYbw/BvS7jP+yJVrs+Rd/47CNb5ctEseP8+oaSFq2SFn/YdhJd5zek+KswtG6Mu91kLmkeA0U
CoB54tEt/N4qGyPsUNB3xm8Vt+CHbaowu2bO5uqWEHQKdLbPDM/vZ3PpmFOQcxDjNrhoz7uGdwhf
KHdKpVdPYvUiQFwKmJlZgpVJlbR9omh9KKJ9QYmNlMcDS7t3uT1o6E4loDcV8j3M4ZqwEWz5svR9
uNQFT1Ze0AvvoYr2gvAPLswxHZXq/xjMcVh2CplC9ucDlJb81+O95ZP1rbrqpp+fvoJIZVauzPeA
iv0bRrpTCy5biGXYuGJk8rmaNPcpPfXOfLuwPIZJMgFIiYUjlvjeUld7days8auSbBQwA/fI0C7t
p7uokf8Vfj8tO9KykIpiG8btAYP9VJDRR3gRRoOu1ainveg/JlLnmDSQ/esPZA+9wdEuPj7rFcx/
/wEAfd0n5aISVYjPP67DBomYEKCxYqNjzag0Z3srQ3kD6/SlVZMInQopItgiqCin2hQDb9XHXnxa
M9K/GZ8YoHcpnbaA0gEIN14fjTzk9qznEcKjOGc4cDG5tJv62LoVzo9KaqnCga5v9KA8LAaRa60f
PKzlEb0ypa3kyZNtelXSxAkT5M0eFD4NRHxNex/Utk/e2apZjZ6P6HLXqWxlRNAHQ6hgWRlofQHd
zaJWOSTUua9Z/orot2t4wYVmckNHWj3aP4K+tgjn07kk8Y9kZWwNRviPZcTkb8ZE+Em3SAbsoQLJ
VP745L1tthMPbvntz5B5ARE5bwhP1dkmkAYFTAwZqW8rAHA+bu7wuX5otyeQdWA6f/C9tPveEYBV
Y5FgQSNb//8g6pFcbP09KbHam4x/yTJDccfe0QO6MWjMoNR9P9UE+4er8ET2NvkfSukhLyXHn3wh
YaLE/UmJY/7kc9VYrpx/eeluKTgJzMQUaPLReXhCD448naSaVlaV7ttsQx6N2wrm1jFhhQZMfq75
APz6Od7i5Lx3eOZxtzyuqCKUDkImHHkMWpFOY3ot5otvuL0fuH4alDp0VgrFWiqcNIOldg7FZJ89
q25mJ8ntGFUYaxQekNq6dzMtopdXT9Cg0A2MpuQU/cu0iLqrTnfSnStOlZjnLlYsO5uSWgZSFyGR
B98utbUZ7lWmtTqXAiMyS2XOq3Cd8Y8rdjUj+RFopowe5s4tMuyJMr25nXJdJHRZxaX3xIy8vVwD
e8N+YcZaDwZDEwyHoELlF46OGxKJM3g+busho+4QVW1BUh0SroozRdtIfDZBFcW43qLWH9iP5AEa
Lg7FLOOOV3DKo0Irel/wLVXs7jDderDVup/JLpfkIcA+ovDbgW+E5CqMTiBvKvzM/fbhqsZEbzOZ
+M4rbf4upNtbTcPjiYxPAZGTRe02Fm1apWBt5zdzqIPBPDAphkSPce1WpESBb0zRGGrgYqwePEBs
aLOSLeBHhQFoBcVBxQbTqe/+1Q12RjDL0PXS0YQpZyo0fq1VrLVOpeGRronEIl3Jd81LwaEqMZce
eEYyhG7Bzhy7G4BPgG3clDcG9oR2Ke1OFNLiSvlhtLNPhZw3fIG+dxavyLY+O5TCBZjuEv3MY8qE
4x51UhtJYo62X+M1hq4ge0BrYY/h25HU4+zbr8LMS1LeBBFhDK7RZsuG8ETjJWz9CcU8XxcR/Is4
EOB9/7U5BZIVg+w4ZNboAAWC9nB7AFwdNA/JAT9wMZRYiQasuJos5lCbDitBHzJ0s5gkwGpMCjJU
dg4nuCoIyhjzOotY55EjTZgCDAtbBRhBWj5l/bC757yDp8J0uJjY7UVLKH0sDIrJRR24I5oFBgFy
1DYMnZKya1kKYs3isIiY4d8ZygLYsfUGbhbfmeS3X6E/jtjQBiLxijexqKaIMgWMBDiLYHlgJN8m
Zv/FZ+JyA01D7ljYD+0U4N3/7FSP7l6MYibj4PJ841pEp5uDM/7uFJ1LjuqSPrNcuxB6VW23tDXr
gNL/DYLTm4Pd1Q4+oK0nn0HyPTUFS1IBSaV6Qxen98Il06yOknpUn+ZNENgvcwfavhO24LTf/3g3
gWoGE1WVYn9mQv6mNGP0qZMOsYyedWpjGGE5pNlv6QMtww9yHJ9mxyNJjSQzB4A2oUiN/FUDfMzl
JXH3w26nK7y5VYCUnKLObkURSE/C5tNhZaiGc6yEYJNqvvlJra9PFOVNxHz4ISi08S5t4LNncisS
CpR8tI81qV54KXFGGmZhn0Ho0Mfc9ifeInq4dhnAMxpkur3cxpHtn1tStfzwGU5P/JQpABq5+Tb3
pEtDeC/xU4XKYtgb77Mby7JPJfzgyonb9LRPtEhhly8fQxsb/pbUzuC0rSLRAltdh2hYvXeAzjh4
nPVyBW52Xuc/uSL9R9P3t0aQtVtapcIaf2Gko/9FAhxF2Y8lG8cAn9kIU3L9jVQvFteGjW8+aJTa
JrnFupKLAf2ea52hj05f+8DGnhxaLJCKYoJ0jU1q1tzf8pycf3We8SvlvqvCmMvqSEJzqDftCdjL
NGgkm8peMKoaf2KNyD3kIzi5IqWdPZC3CkTEu+tlg8hec5Cwz5tn1vPSkxsMUlQbxXBGckfYvVed
Fv0uMCdekrIk80S+yGPPL+4ZambxNLXKEgqIMn8V6nwSyk79omEh4Y7LjjpmN+Gumm6xfO9xrj4g
KFOQ1zzpOOJowfA/5i+CKVVlEe44v0UQio46R1kE4bvmXySQiN5q+8PdLfmw8DyAAAFT5b4U3r1B
iFbiHpouWIfVzeojw7VT2m8w9waEXwOSKmIm1XK4y5qjgDSQJNI7/E3O8DCYIks3gfq5w/MgLYKJ
x/XFaJha4mmVzzTZCbGvyxWk48uThguoULVxNgeVFo+wjAHFmIv3jNKhn+RTP8aJKPbZp8Tv5oqZ
EsY9Pm0vJdFYFk8ENvHnaA3jkov5B3BwtoJBOxj1l8hec2lGh9i8Qi9NaH4GBW3qSrmBH3oDB0g/
tgQsSpdwEGQinv3NzsUUXYaD8vNyCjTxwMpa398H4hrMImYk3vUA3CbbZvc1HYz4z73+ME+aNiFo
tP8SENBi0wL/bOdiUjcP71wb1eel78UKIgBmtnyYlM3tLdCJO5rRdIG32XaiuJ1D4/ZR63aAPrcV
480WnnKmIdv7qtvkUC7Nih5HjBYkgWy2xexYxBflUtSM0SlroDfFq4VVcKL+7ntPh2mH6e2ABhjE
g2r+vmySAQCXJGFaJyuSYyEGm5p38e2bl3G9p5jgZ1bxwq9DZm5oUPfGNRlgqJYQfFz2UL+kt1ZF
XS5iqidS/5Qvnl4OFbiX4oGjLn+R8tbkEJ/OnRMSET7lOWhvNDCYyypkU4VGJgHePwsnb6bLC49E
QkmLFY9Hbshu7GtCPcw+1gMcpklMt54E0NEDwh8oHuGi2lyGDjcN/fKeNaMctjeS0VhEsGzk3zXZ
3MN1pAurCJNRG3UFt+O9lQ3NBzlis5+nuiOSoV8H2X4pOdIh3EUlognKrPPfCPt3NV+gsVRnd0YL
oFLzkKXKDVMgLNjHWYbhMYpzkhkcjO8W6o9Ch6zTmR/MHI1MCpQ2cOpfhxoSkd0PVnk6txe2SD81
yvMaWxMZVOyOThIx0bJEvM73bXEC/qJV6bw8AjRUMfAjbpdQByeE0AbuBXMSKTmcgG0FDnw7K9xM
VRHRWbAUgW3kSFP8DJ44yI9SkxyT5nBpRdVgLBVJVLVT/DRp6dhZpc//2jzPPW3qxVV2BDBpwgyg
BHhqINSzFeseG2EU9FuAf54rlqvP/lyDxGnurhHeEcsCcDN4xQiUFz6vFZKq6jISfKOmaJDciKn0
xIAZaZdkkmHrqirvvkPGBwukrpTeMsgi1oyVZuebvcTcpZzSHkwGSI/y4nb2/jrZ5DSSqGYXpSM0
VSuhN6W7yvKqgLBhZ9LfeoPmEXleA5iv1hcMSde4Caa+a3wonC6DO7CRPDGA3731JZlRH8krgRdY
UO+/cHJXfqTuizMxAQKvPEEwdacbsflgp7Kb97PRtOpklzAKbJ4CbuDEcGuZXsjrp/kfQjFHYfMo
mpgtOyD8EQYa6500mlv8JQq+14XqbmPGPqoDy5zXyBjasNKjI4fU3gyVCc171fmX7Zui1rCpSSDj
jepN7baCSx+Q/2KE/jXN5g/0VQI9jyb19ccUjKVN1Md38MdrQkX2S2AsiG3LveGdGkFFQTORwJMD
5dzDGL/AxQte3PQPDyWjHy7IbSaCDn9KZO+Fk6hlHrF+OcG4UtMlK4CXQIaaUieXWYyjEaJH+8+j
UXSEU5+1SYmD3K1h2+4kFIvz4Fz1gop3jkUQZJQ6HdDrmCag/aKd+KEtutrmokcpzhFYWE7K1t9B
t3rbyArjhvJx5dOs+ZpdVVUS/UU81GPz3RdaogpxFrjh6zqofUftDwroFNFr7SyzMuYH8o41+T0T
e10E+H1/tr8D5bDfXj+qvX62f9YLUYyb04cb0IvAZZxTJ1/g5zCJVuuc7wxbRwwENGeMhsNfDBhg
yfrwB/GVQy43RIDk3SWVNObGpXa0AfW+xwLrlVxYFJns2ZxNLd3BGvIAznHSZ0RcYFMuZAp3wJHs
6BtQk4gwjvvS70bu7kel+qqPZsDx0DZ5n5ToL6lyb68yyKBOM5QH/KUXdz0FQqePavL/+hrG2F7d
yrbvuTiKWOm/yJ2Fof2XwoZy0pJVZxHXKvJHi8NUf24jxO5ImmZpE+ppZeEpa9ZMckKqRhVnctnm
NCSG5W04PgdJsoQkOuXJSm5r2LAgTjD5Cy5ALH0WXr0KamAly5NJCIqFN6azMWcNmXy9/RTSh2L2
JSJ3Fq/GciQntqz/r0KMwvOH50zIluo729u9iKGOuEqtH7P7RC7KtOFbxalq2sytrhpbLjuCV2N+
Gd5uTMhnaodcN7dHU4VV9qXWK/DO/sgIpAT5Ku9tf8+U4JFlsTEXUecioWdC5xKYVJXQTVZqEFlo
AF+L8m6/VFHfumfk6PSIg5e8tnzJYYt0BT8hWf/LjYsy3BRPU8rHZvUa+4SFM1Qygf+3cz5kTlYx
TThnbJWNl4zSC39Wd/u+J6IEMcZYgaSNgo08B1H9OimEpj2Uzw6YeyVymDMX6T4a5vrkBO5EayfX
0P41D9Z24fa+bKAblCIc3SF+4rcnwO76CP5m6AIV4oXNkLbLRce+zyr539gRTqHW3oFjKwj/io6F
lS5UciUeeHV4yrt0cP3NVAR/q4lhGLFvawi+o2kyIN1YSitzej9UdJ3cvOadfZiqHzbQrKYFtqos
h6ik7KIcBNScLoS3yT5B8aADf7o78ugpYrcJEalVjHfzgNVTYruHkLZHFdNhDMfx/bWOGbhPGAGj
jCxznMXPtR2IOm6SLQbUELfqfvwRohOFu9kkq76LsC6ku/MTCCx2sqdxL2FrwoP+GbYNCui//gc/
RM2HNoj5HLEP490gNTFItZtaDtJchIIxQMKfZ40kqWCr3MotbtLWIN2RneEtz6dQZA3jD27UF7YG
ofrKR9kjvztCmtpuveEw9fxktRwnPYcQmhAsmyfZaIkDt2M79V9LQC5ef9r6OPq07QIGLoM2N7Tf
FyJbOJ2VMcexayn+lHmo+uvI8nB3BcPsevdT73noyhAH/bNM2/uIfhErIYxlVLZ4XZURkDDsC2wq
Pp45bhKUMYbkvz/ozLePfeJ5EPPtpvzUKGshrkpUHyiSbPPnOznN6HXsmCNQDs+t+FU5+4Rez3mh
d3857SdOPNcRtT3vuLkLz78peRib7htCrnGmaAl473f/uTfk3uaSr0G1qP2nhL0ZytX9sLoL2Nju
74J/TK0aZYJaQodc3WttMfWkg0ay/VKuBHUImMp1wHdgR4MovJ9jDVAOtMkm7NZDE0xeieH5/8VZ
o6PkB3t7TKZJ3uII8NOXnMi+TwvfPt+xkaQLMWcyJswxHaSX/9m6MS9j78mcaUpuHecMxzDbBumv
nwKLeOLiC2DdO25SdcFH/NWX4cMswy95OxZkw41PNAfDQ/NAr92F9CsdLfC0svOdAxo/qJdGeO0t
WW1P8CnbO+lTyGHlBMtJ9xXya2nhNzN7bjjx7i8zJ4mG7pIdaR6fgn0eg9C8TJQ+qDsskgEBy9tN
V0enBzZNziNIodw5Lus7/imU6tFsif1vJLjyIrpVwELcsMhVQAgR0nmEBKWDrRHHF1Jrmapw3TGK
e1WG8i0fQoAwqb2Y7jYvhKXcYTs9BmMb90Gy653xgI/35hSPXUoYnb6wpK140MiF1+RHL7AX00zF
wQFRWFiZXT6bzcBTcDnBCi5T443NwH2Z8GU151d9xOWx/vszah1jtCOd3/GEPCUHgarPSPB1hE4Q
jmftNeud7ukQqoOVgZZ5Q2IHl2sKl+94sd9RUyw/HYk7itF/ppdLSw08BK1prRKO4Kuu7zcKMxIO
0MQL70mxdGh2TfjZiaOZU082D4b3qi7yk4YMcW2DCNbvOgVZkTH4TCOND/1VgIzyLwUl55nhld5g
erkdN4s3aVBFpNFIic3vB+BCheYmXnfbgwu+kXek0qZ7D7WzNZPkRcX4ITBo5sigQEze4CPHWUZ9
DkAx6mA/OpVdFBmRDscRJy9nYCdbIH6fK0stQW1h11kD0uCeo7VbplEuHPkrAVJmMdLa71ImgxNu
i9hHf1fiQW4DGoSO7hH3w/uJyZaJPC/IbGb6sxr9vBVDVFqqGFzUClKXSwI9+jLhygAoqmWqUXEV
rYAU2Gq9oXaQ2oz9GmGuh3VnUZAIunyqOcA46mw6deLgAimBDrRIUpV/48z35yKUhPU0r7hH1gTI
aroYNbVA/rXWEesQFzSvvcnzclCRFe+XHKoHySbhkYrqSHSRrtIwzns0K+EWUw6EQEKTxP5At/1D
8n9W/DOD+jT4ZFOdUFxYzZZd3onUcddtzWMZ6cEnuLQQna4bZXRTddxl1GTUHiir8eHNRktQUi9/
Q+AKbq90AMkBTk/D8+NcT2sexMMENlN1A1xLH3af5nHXxRXZys5zFM89fxdcZqzXcVgXA7E16P9S
d/tMWVNM2keRSMKnhu3XBnZyrCu3a9iFBJztzyPUXl5ZVb+e5Gs9MezJdNyKDuPWb7ZK7+tXae6k
3qtHJs/M7XTZpVY0DlpAehtiJrVOrd1bfxPvH7xec4QhOWVYqizp2eeib+i1THW4nVBK3QWatVyJ
FNJzzB/GeoxcAnny4Edfyf0a+d1ScULlEVyy1sMLlZAG/iZLl8fb9vRC1VNfgJ+OXKYnBaXHwyO5
noRCAEVKXWlQ58C9JHBgWv40FjHXwm7lR+x7MgsbHSFHdOa4Kc117stsKexpl1DQCiCrwpu2bS5A
0JnDN680GAoPy8+Iucn55QTgUADAaBbTy6EE99IW3ZMl44vc1zPdl5QHQCshnbOYtSL25C4W1R3A
/nHp91qCy+8FDdG5TRVr6qy7qFlwlPiwyhm5ZhjZeK7ZuuE2RdU5be67Y2n/DPkUVOuiKhSsRR62
NYO1zU/KiybgJ1xNF1Rk8ZWFEQnXdW6ifmqRUeCdbC6z5b3/vWL4chzaSy93MUvhM3fuzOw9KLob
5wx9M4F42VS1xgVX71NsPC55FLmqYe6mL24MmwYZaXELGom0z+mRQMDQsN88+L8xagB476AnwtAi
LEZacP+yXeefSAAS404iVwavcUmOIjaSNjuwhVfS29icL71EAmGE6/YB4lwEY9nMkz7bwpOHHVXy
1aFlB2FVHSBAw3n+ncnJsMkfXMEyMFg4LrjsmrDeHk59SBtq/zsZluKEDVSeo4riOzmX78TMr2XL
C5z5r3GrmbdiU1Gl86NvkJk7iXYwJcIV32XNycn8cN9k4UFK25C6nnYDq9D++cFIoWeSSn5A5G9D
56Zhk3I0RtQuFDkw//KF6r1n/wwte/KED6c4AeRUJtzmYXOFKa6Gy621ydrgM/m9aTxmeD+9M1KM
KwRVRZCcnYd4Lckt28h1Ce3B9nZiXW/6OrRBRY2lV6+fUEp9xEeCv0BsAh4pWQ3gDYSJo9OwvfNP
qzsr3/C5cdhZC33+w+Eo7WMquByIekAj5Swgit6PPNlI3nRiBs6+66q97p1Kv43Q3Zj5h+eRP+ag
afOQRIOd/njGsNnA90zhAipG1SevFP09QMM0jdc0a00z360mxSJhnGwAmQlb8lFjoov0MB8evx46
bORZk+crAagU5aHs3KX85tPVk0uoWBYppIwNbmvrU9V+eCeAaBYaQ2Tij91Ts/NhRm96L1PNTTmj
f7K1lkBfJim+yMl1C8tvfmp073h+DlEYqIRs8q7+mv/UsrwVTSFOt8UHstFzW5rkZNK1/flWhAnS
0/UnCrNUGLaIPhF5dwWEWI2y5ddcHapghzvSlrSypD0zZuVvRB1r7sjT6lZg3oPldPJTjUmXhKdL
EiH256q7dacSOHXid5JHmwiCJxzS8mfZhd0gB/xCJewJDhCcJReotcrDzD4NEE6y2mIXMajr1d5z
a6PYMaGBlrrd2gFk6P48k3u3LouRuJRk8qoKB2CyM7s75lC9wXWdEA7NTkIhA6akXQ7ZKMZU8yDL
M6mtrkGcXdbYlr15NU1x21lwfqHOdFJgYuAl3aVLkZc6YMNUSvYmXdUV2oK8fX6MQzpkV8YVCR0a
HT3/fzOQIASQQ3wNuE/fjr9kBaXSOleXOGwwhsC8RvYRGGkIolRvzCJ+RXUTPsEcdJa5jhW0Zn5R
1pxNMZlQbM7nF34g5yxnYMVmp4Um+d+JNWrSS4O7l+qRgy48BD2PuUV7Uv9J77JsNUK4uK25fP9z
OUhRQlJlpECQsUzhKTCD3rPBgXgoqmW2/tVkS3g+Ke4qteP9iXxS6akFJXgDXCnWm/HsU77XXtny
JVWCjktuwCYK/pqLisXviXlmK9j1yyc0Y1zGdkoo5aInKduRSQASS7UCMoTWX4sIRRJCWFIe9SAg
tUwczwyALllgP34adwpRXwucQjCat5BYcyAO59qJ4pI44VXxRjyIeHgLeYLdNzHvqdIIJ5mbqlle
HmwGEHlAmA2O06NS3SWLxmzfmnVmi8kFVMTxObN3kfWbB2/S8nRc2VUxy+gZA0izCe1q2Y603Huy
wQW/OWoxXnwa22+vNyMjMToq4YNDCZiU4COrjDGj7wNhQH6OIlWQ+/gkKReiMiZVaJ6WaElSo50N
QwH5wSAp4Slquhc7ouO/S8MKr3gEw7vINCva6sZCziZzvtLSdzxoBzD6fgfQJxfsfKOGfexxEr0I
f9/18CIjCz8MWIV6xz+CcLDRblEzHIZSrDYgjxaIj0py5Be2ZtqDJVC/zVhtp7PhNN+jKSWsY4M0
XD4oV5k9VO+hGlV6NJ/HFMAfSnUqIpxp6An3RM0ozjP0A0MsNfqgy9U0D8z2NKdKzrzYyfVvYIgw
Qk8LweVnB5PSECBuCfA/lDcIysEfRkwnS2O09bFMkBXGLpZv6PfTFLd7HZjRPO230oRLqPt2F0IU
yFZHTixkU+XJ2Yzxg3z+6OIjhv3dIw3gFmaYp7ul5aWlliDj2uCK+J4kZAxE+/sLKVi/ANsAp5U9
Jz9hDLCWY+FwcNU7b6lx/qOe93SPXYcHVKtOrjDDxvv0t6109DcNr1kUkKJ80me6J4lvztvlSWg4
/wlKaWx7jxj2X3wnJ+17ri8gtEsMJl9vL6TfqaSY4Yg3IhvEI1vNkFPPachb5OoQ8fZaOJmC+9aV
owP0wRz1YXFKNg4Kt4Qh7IZK9mmSc4/D0Kmi8jW+EaX+3hXo3ru0rwr5NDoH4y+/T47UcsoceAtP
KUi8F//RjA6OyMEwt3/uU0aar3iQbw+GkluU5yD22PT/xaIyHIKf+RVEFA4XKV3/XqAup7eE3Zte
0k4BFwVZiS3Dj26MQM1SEJFmhyrmIP2Kp48JOYS+XN8Bx0rugHY/VOSw5vfpKgeUnHFg+SIIpDxp
pASnlLhUS67EY/Oklqbrh6FyLtb+Cp/lbmi+PlRZJPCeDCAcnKv6IikzWcxe/YmzHUfBpcVVMsyX
FpzKv4Xy1k1aUp/aGhzAqKc3ybBjxPp559YoOPPBzks/RoEeI3cbosV7L83ka8SagkS7vt2jeUNF
xxgtbKo9syvEDXT5+CKr3GM+Z9EH8okDB8qbrW7tFCla5Pb8rih4EeKoKzmlTTvSmYhlfyyM7PRE
SjLiD2Mzqyd/ULxc6RqPXb7J5vd1O/WtUmy+5npZ7AmBVKsHd6QTrkTIm+9BvB7lxdtCRe7SJ+2S
iV72xIn/ykwVBGizhAnzjoVvENESkuO7vSBH/MGy4E4pQHytu5XW7SafhsUM4rrZYMH8WktRV669
HEJ4eAttWSAwBCA8UdaHKvMatiXvuTdcvL/oktF/Q73SK+BMRtI4KWqUXFTM0kcxICxaXYdLO2ue
VigI7AjAZy2k+YU6tklMyG1vJUPL1YxgbzhKKmly3Mw7tV5HZ+WsuuRDcoMOFpkFLmNsA5ldWH+F
WtWkUaWTdoyVrva4BQt8gfmsrjpPReM2SY9xQBi8ouDV4Xbd+8//tWl9ApzXs23xy4OeqXZThhgD
NmvH0vPzLx0HzUOvTwoVcKByPHBw8+zhwh/1wkjPLyeZrs2qrnw2qGGYZn33mArvIqbAw/Y5Tgi4
knY6d+ua/52zsYKOFnOXvyhRuTRCihiudwbnvgvlRoI5cZOg4IPrKgUauFDN9B/XzHtFN4OowIKl
wmXtiMhsbjon+D/U4Vu38xyoQYw7F9p11YktY3g2amwhRDgTz6s5rAb2UP22f639Y4x8edHgIDX4
WRmf60JXnPp3X/mEPiWeJwjagjAv7N0A+H6+l2OtvMpJieLdFl3oZnfuz4P4Ojr+J8hPOrlJI/6t
ANP7T3jo/uqdHL4hXqb/DhSSLE+dOqTXc8+qBbNT/vAQ1spQq810eteM7Vq2cisbRnBEIpFGwBQ2
IBY3C/dZelv/jKPN0+oZNQ14pwCAILCNmeMjeo08B/vr+tSofXK4OmU78N8deawqRNlCY7I1UMWr
R6HPsIaJpFsucYDdPjdiNULS56UT48sm5T3KzCh11BIvErzi4s3TmFd1YHjyHdAJc5jSe4zmiQNa
gyCa5JW2h3pcQO1f4bBnMByMH8BZ12IohgdIBTp1E7DG1o/7k97+uNtR9ENgd83MfujWPsG4we4j
Yi/C5Hr04ttUzf3NsOW1B//Bbpm9IWRh1MD/wrjE+Dk7F4V8Jb3DWJd18Sg0uq7KSblQwZy5MQSx
tt9Z8vohp34m5JOG901FCnPbC8wp4QMsQH+3/7rJFnmXVwJtrQsTblW/So6Xjj3/pup6m0rduLaT
aoj5vMuJcKEuY6uNTVmxRMjhiRHpCwFkrIhrmAJzqg59zFROvwo33sar8qsUaZL46rXNjU4aJLdx
XQulZV5NwEGdJJYR2s7EUPXf5wN/LO+8CQhY5FENV+BH9LdU9Nu+NgnCi+XgOaPcTDzk5aO8sp/I
VtW8XDPDN5mv/a6s+AIeaKVfW9lUjlSBBcgRUejFRqh19uEwRTliO8ZmK4+5lpt/e8zj5qpPhs4r
46C2QabNXHWxvxvz0A5Ph8Alf+Ua3bl5JHBSVL6+zENip+6TRNCytV8/fzwrsHc8SokwioBzvJ1s
HB3HNIexo8dODxDFrhK9Pd/PM6l955GIAsjCaU6H/h+URHT2nlfAJ+PhhACu3TpcwGDUO9dvT5Q2
at8LeWZC+3ffvMea9q46jZ7EdHxnDum1YEIZQ97TKhtz9ZcxyY8DS24qjXIwaseq1M13UqgvotpV
U4dg15HF27rt0hS0zFxwWh2Xhf5UQQtG6c89DreV9zl+neDvEMyqI62Nn/UG9dry2/QUrzBuP79n
scfnpSn+uOULGrliEdNx9DbXGeCQb+TQaGKnIhtr55Zes6XrNKwXca25zMC2+/MLrWyPZQB6y99j
/DnPZ+vFpd0JbO27iOT+ZIzHwzZK4dfstODcolln/DUFnbQGvzvCox/sE2ZPJQa0XblnpRk3VcFs
qLs+mzYzSaTX7wFeJztQsz5h5JWBzAaWUGZLQ8fuknp/dWde0rVI2LmzxcgqbQk0N9EWty1MIUcS
/o8prIDHlwL2Jw3xl3na0dhChlZjus0fVyecUJ34cCHYDsdlzVMhwGNvGkFCocHY+grnMSl7Vuil
HIhtoX/Z6Dencl6ekvrHko/Gq6m6x0laJOlNfQLs2XXdnub/GTsG2eU7JUauMtspqq92NA1U3uKH
TI2jJ0f3Xa/EUnDgO9N9MgwgSKu+eJkozuv8UqGsS2D9kMoV2aqaDuyRhc543u5e5takpM5ldu7F
7wozD0qnYl3MQLwDwLkpZnM+SrHQ6z56RlAyXe5HLYK8VLbORnVYuqou/LtuUyiUSJnNl2ljpJ7u
Raa0Byf/216MFI16mXJBa0e/FFXz8CIEarlolQWO01XOocHmoM/UNvU8uZVadl7K8vDS1xgfe7Wu
tWZYRzWOIElf5KftaKR47TbXKOMQ1ez8aAj7hkBmjayIAUjOJlpXVu8JNVqEX7OGC3xEw1xH0Vyr
f124VflFm5gZQtFHcU6lSaU8usOdClSvwPUVi0DTZeBQhnW8ZBOHj3HlYtQaSr30cEvwOC+YHYh5
WhkkZcU9bv3ER0MyOrDj5OE4V4SAnE5c5tXC+OpEhXaVQ2eL9WE1ZqA9lfYsOgeFNwD5ka4yG5o7
BSGZ2ebZG2dnlZg3aBSWoNRpN0bF6GVj2WHKYsBkeb+Gleamq/8GKhQTVZAOu9rp2RrDJStq961r
WqvFjtJ3uqRlLdv0bu46CwE/A18Gz5lVZLQyCIr/qwrwoUkU46cJ5yY1wg6UMBL8C6bq9oXzSyac
OqIglRY2INJ2V3nJ59CTywwbOWeGOKyq/plcvIOSOnUJDXP4e8bFDXIRYKHEzSw6xYW1zRdu6OWc
ukQwXhZCedgdSZiSy0ZVk0nZSbfuAj5yXwR/sEdSJTfUEi5cDhfSyaaC2I8Q3dii1/YpcGxj/Z4m
IeGWKUSf0xXbIFH6fnmnX+K5bl8vCdGMy8AmZ692ZljoHjZVxgv+PmzuoddnGxSVwPjNdQfd9cZm
eN0LONEy0X3Thzin3s7UH12ur6N7LCryEVHygDIXAfcI/MwXXNvH4ns5gEcCkwL6L+mm6CEKY6rp
GGdLeT35LDqZd7QNuPAjxblbj8WePdMl//e9Ag4ghH+zdbfj2XdzkJejnoVnLIZHr9IHi4Gl3JcX
mcFVWIuH2HKQesEgPxqIxadbJyqFGGrdkSd5XME9Uo++NAqAoN1/aow7J73GbFLiifNLw5owQpBi
uH/xy4mpGroxSc7EQ4Ltuuf3SImfdA6Mjtq2jYNbS50X3YdqXnGZfwxiUVY1Eicalt2ewBtpvjjz
5NTZL4nw1Ci+mFYfsk9ro61cXW2LBlXS4jqoXcRpyfm7MNJoUS66BLuMrGm09ING0WVvI5BrMn9s
O/nLTh+OOqXBwXh5Xl82bn20b9abCv96Qb+PGIpAuJF0w4GmxsjR4PASkfMH69V5VDRX8HwNum9N
FrCacno7A7/fMWZIeOzZP7uxHefI5AIduSAh7JwngGROCPfxrf7/GzRL+MAwOR+ST6NnTR2hPTVm
ClEnmGwsQTsWdEbL+Ifaaxv0i6tp4r1hl+boem7AkzJwEjR8T3E8YRIVyD29xcYxUOd4gyImwvax
fzhp1tmdhSiBlj43T9tEHUIPb1kThLiGnfNSyuIH3HRLva4eq9Z6ucKJwivQ/S62C9mDKyL8hm2B
RcdtO1lHz/1wEojcE1fYx8fnGdQNfTUSbW/FObwizR1lPTdyCuyXdwtuPezlR2SrV3O9QNpL/EmP
f0calVZi6v3b61n9vncKwisB4B3QeucdO4gdJKrodvTYpUIyT0U+PbOYXtvMp8M5A/q8UONSu86j
FE5mdyBtxsxy4f6olpwAtOxN5jWFbX3b9QabntraYjT7EOHowdp+Rmzs5pqc0KaGv74I3NdCzJ3Q
TI1UzRSC1ZT51J8ET1UYDnkpClinZaNmKL5KNyfD8GqWxmhElS2QyvH1Xq4pUh9RQsqdHtVzBdqy
rHUx16mgvwXRptibpMMlLoMIt4pJSPf0K3oEGRMTNnp3JNR5y9k/jlIBOVyeyyoPtTTBXoplrWOt
EtNY/3PU5p+8yRAy9bkMY1lbOWpwQQclXJVLQqUcM3wpeA597DSW5wDmGBCdPWNtQQifocoDoNv0
vmMvShicjcxmFT64yOA7SjMudIvgAIYB7nMk2y/linhVOzQt6c26r/LYZxC8HjSqFh/ieSodwVjT
fKFWukx7wpC2yr27EDxXvvsi6H15kMAD/HsSTfoUoW/Jz08HmmnzLY8xmZjNop2GV+Y/4M0fNqnX
AboVlfavJUAf1fZifdqkUD5ToecowEE+kmPjlwM9inkKx28e44c0ujsfq7h1UIOg/9ODrOTtnQZF
TassgieYF2gIBi46jytvL1FC0/jmyofKq2tF2icEE1MYyZUIiXOCKtjbsKEy9hwrPabVTPCPm9XJ
1Uay2QbimflNXPWwpGnbLtUCxup8e10KTVH0mqt5Pz/BsYF679csGbEorriTtg7wbimEYOQH4Va0
yyE2sZvXLRL4G6aao289v4yz//CBlPVXmmNCslac1QrrObvqPdKXzdHlIw0Zid/HDOht/xtWAgGi
VkiagxQUQn9xrzS3mM3wd6YpbWkkKNOGuvxM5Mb8w6+nlKU3YilUZFxL0FhZ6oYx967NXNFdCNK0
YyT5wVPGR0MQAQ1EUf9KSfzPryNghvOdDF0LmBQVKIchXFwLvaSDLpU/GFXHfs4++XZtWwK5wdMN
BihzGCgHgHAO7S2AM3NOHg2nuDcUp5mvgoPyEz+jn4unKgbcaZb00EH5gYEkZslUgQ+k71KV/X7F
w9ShsQmFNqG3MDpNWladU5yMWrXonPGqUSR/GBb4R1/SGjWdkGvRhl8K8/qNtMI+1xw8n4gBUVd4
NGX8lWE6490pH9BRexTS+iREesRGpuOjupD4O8NbrkVStM7zkJQwoH2stIBzPIpte2rVl/BTXPm5
pSRomXkfSvHv/pZ2RDPw4YxbmR7WI36o8kKvaxHDGNcoe1zzLpAdDwWMTmPDJhZD9O6ktSBL0QyC
O0y9oBGAgBwL0PGNsNYxhQE+Ui4dzJOIK0ip7zuiWRrqj7x0QyBF7R6ZhkuJDrXnc2Z88AWtEDSn
MJTAF955kgtwy2s3SWVSZR7+dGHznSoIi9sBbpbY3eijdTOm9h/VGu1Z2jL3CyNGXTgAUlk0evs0
ufZ5U7aDNIQmAbKR0Ut35qG/AzluWeLRUl6+L/wqwryVIm9+NUMLs6HEQ0PZSpJYSS6U3+0eIWSV
lw+9Zt+ieqpsAwDjON4oxJ/f7Q+cPr2wjYoEI/OrYpgsJMj2M5eC1B9XGdfACdH/VcN5jdV8A1UN
9NCvmai1XGNRozTirnOS3hSpvKSGekbeFWCOfvxhRluczrpxKNYpGpgkJW82QHz8OnBz+dHzkUaC
iclWrOKdtwIWDIr+BSgjV0GxgMdKyC/0E5Ue/12GKM0si+si56v5LFJrGwPCGJiKKnmcjOtKaDtG
EQT3R+DNvR6bztv64/USgEipZQbE6aRGlQYY13rIrK7QvGR3tbNyFLZaYUoNeYvUi3jD73FgQD2g
tyIhsz2gu40f8NEmnkJN1gAob6rElhk40NybJwSoYgMQwzI11wD1/7o30Wfg7Us9MLLHrAQBC9tY
Xgn/e63z2knnqoyp53+H6uxp4QcnmzFhYfsxNArmTajl8xOmCQUP4OlS8fo3/uwvkGEGp37r68p6
THJYuU4//l1Sf16nY8QFKZ2Q47/+C0NtmGFfO0MnzoEu+WId9OOYVOpG56HIqMffiiMKu8xtx5OW
XdoChTm58wFrUFln/oVeQvGiIH8aV57ubIzVanTl7LtR/eOL/x+QlFR/rmcDbT42o3gxPuJdjkw/
st01CdA7UWp1GP68BBFsX81VSwjM2SwToMAfjqHbPvUF4F5ghTSyh2fiSpJRfoR7bUvG8o9295Oo
RHzsunRGL7MzxE+uPnQwtdkke1pCfUl7EldLCjFHh8VC8Cy8d3ck5Dt7ulvAWmcg+997CDCHp0/W
Z7/rPDjPmk5r58fu+inmnlaQKRlQKXNuXf1+kDAqVV6TVOt687/DAcHztr8FVYkMEPvB0bAGTXIf
xc6t6R0ADKjD34cUkoCS8NbIQ+NPXFMgt5UfVuyZcy2XE/Gvg0JymJ8YxGmZyUtm+SxeyB5OF/4o
K3JGJkusWf9U2UM62yI4BQffWTfDb578oXwN+zTRpBkLLWrVqkLvSkSmB3T5hB7oIjNMQ+XNC7JT
nAgKU/12FnSSlST+IDMUYzXdmDSDSWVuzms73zvb4kCatYfbZ4SM0NFw+/63CjGbxjQQsNGMKs0i
/9u+Sp97WOBXpzNXwkiEC4MfYYLXdGr9rp70nZk2Z8RoX1MeCrqfu1gGuG3RuRE9oCDgxr4XiR7R
pTYRQSMo1AcQa9l3vzrjKCTUV0NgWmkI63WuhzO+18pmW3AGtKc1r6FfxWWiITCr2LolLp9UAZH/
8cyAGu5wN09L6vcXXmkepnxQrxzuogzjiqTu2xGrnecvgIiSzW08YpFTuVLjVbIOgn7hHtZzVP1M
nUlNZCcaz1vS4xkbgMET38xynrpLQADt5yyR5AoWOt7b5FKPwBcfGQ2vMH2Eu+buwtPss9b6tdV4
v3SqNZ+bxgS/7/dDJTWmERUPyNbwt8Q90XzQy2HydlBkhyqupwCn/RneDsrvWMC6EKuaKkYd4qFW
9oBHuphSYclZhUEzKLJWXAT+4hR34aZ6C9x2zOimWffggkNsJUDvZWo/K6T1A7600DtPyzQ31frl
DBhd6KOND0Hs388EMUP26gM6tbiySAaVtAukDsX12zMABSZzer+pHQaUPZ0Mx0DiuPYdeYROZEWE
VhRmdOs/BvL8VjiEOSo0CQzLXE01kKvBlb+fi0Vg3lFv4j4rCzVCG+ak1Ed7vHL8rGJOpCXMbjx9
GFF0UPKTpx38TGHnIJ8dxQaUChchjfQ2X2t8KAhhUq4e6V9Z93flYJJ1vWuoeWmSy8uI6bkjSkJp
uJEiOx++VeFoGFryUYMXsGRdOak3VlfvH2ExHWXM3Q3NxMAayL5pb+8+TrTijNKK1LFZGgn0CM9L
O5le8ppk2hiymhSqAc4m/v/EJkH0eJfBNr+1cy+NnYbEDDuFzJpf00vI193SGwZWhIRrq0Yw0u+3
Dpm7PC5E/ijxQ45Qp4CBx4ZYcIIguFNgak5gFCB44kmwCRHwyLOEDU7aeCeTMd2dBO1ET2yWgqTQ
TUmVdEnJKZmqf1tEnf9kzGX2PPYO4tZ4I0BsvmMVu/538uUz04B3Lj7a6gGKakjQEsM1BDfrMWNM
9O0jYHLi4Kkz3ze99QpuRaUHX1dDFcJIUT3Z6VI7c9IkxweDSlQnv9wz4yCCTChmzlkpfcS6nXGW
TrHOjF73SOL8AGfjOHuWX0CO6Qye155xF8huaUhhdakbnxatgLMv/9o5wGOt9U/i5Eqr3Xpa2F3z
aEFELcA03gQvYJnuMlO7cBIWaI6LS3NvNv5W7lX4L5W0szVEXxwFgv8XOB4RqMYtBNNlZdaNZ63e
Ue/jvzcwhHsH86B1t47lPj/xgrGyxlDX5BJ5+ir2aSFr+n7nxUIGQjbHpz3EkUqR1LwDTcicHrhS
pvl9N/LvmKSFCO/y7gqhYlHmsmPGEr7kHYcgTw1t480Qjt1DSwF/lelctskJs51kr9Uk9S4I4/dG
wIf8rVrWSoISfkXffOFYGcC+C+k8TLwi9/oc43mIVDFM3ctw5kfQsi2YObvji4vBI3eKPEuddWOz
/BhvIJ7Oz3tik7yUfxp2Lkv5STRlyJoGoE9PFVQrhb2qzhLGwX0hahbEw2FKNFWPR3bTpd5JUp1u
995ZF9sX2UhPj1gklhr1U9oy45BODXHiqR398izZwMipnqAM5H7O83frHABepo1IVeOKABhw8dpr
v5fm1sxd+syL2r10/7xEZmT6ltpWOzAfH4JZX0kd6yxkUxEIQR4W+ohRJz71GUcyjq8CLbBVXYCV
2G5YKKAyLW5C2cnCzx+FDrXjOzky1JsnEWLvrkAZUwNKQOr0r+RlRIldTzWFmsW+3Tlsk1m6sm4p
QAhyUJ88Ki6No/NWp30RTGaeQuG69X1LhTRscg+PqWshyHsjjeXbM+lP+yWu6Z/SGaAFKmrHdrRo
9Efuk7sd1JvqpXcxdee1mWwdFdpO1dLEF1CzjdhwiCvE9YI6XUmS/TPjiMR8IcrBz7hjBbn3wKq5
/144UNfyUHI4dR1eBJtoNL1z6Cx3CmkUbCz3FZwMFLcO08snJQSwtmE1PA41vObiZNgWOiSYzIfe
mlvn664hn/gF/2SF/Hb5sLO9dDREInkNF5pBQgwNswvfVuIperyOQ8vzS8uTmJebwRhKd/et0MHz
lt+Lc/6eslpu3IYz85BUVON6cnqH/rrBejOEbz6bQfgeJo1Qp5hzAfABU1znFNOVl3i5KWkwAiur
GXTLgmtJbJ/QsLSbOkAWFlaReao2kpwaomgNugkM9VRSQofeEjOef67uCfmG//enV/pswZjj/T36
46t0r8nFQq7dLDVJwsEnlJnuo1TokJlTAIkpc5juH6dZbx4KBriO4a+fNQieEWOfDW6VXLCGXbwy
He97ooTdD5S5CI6MmPYQufiI7Xg5aN0xUjL+4GkevR759AQaUdJx4VIlBtCMWq+bPZNMdFJff75Q
YfRgBb3o+TmrvvD/IdLi4isyvIh0Mxh31cVG8N81+rHOSmjvXnCe50wzRCFa9d620wYdaSdsXoBO
kcWc8KHede0mHxVdA1ZxuRlCrnxHpFO59R2sOZo3z2HY/CFWAXFLHZlHpc1z2Hq0q7ASgs2jxGC9
3qJ53DNsUtH40QnxGnPnr3BED01zJijQBE9LbjGdZFk2HpysmQEwmVXvfuJgaIYLjeFKUkfPxtd9
nmRvfXB7B/RQ7J5ALT3jImoqkbyA2OvoDQ29vOO4veXYdrtdoAZoUKJYPx10i3HrKmiMDUUKR9uj
Si3WQzoD0dz5Gv5tzaJzJk92XjHRx9uP6v73p5ewnBAWnJ2DdlnkHONIRc9ebeTQQWtndyVTQtJ0
z8jqfbNPlwHEpRJwW+nVKDzurbMzQG6xdtBC7Mjq0QFGdVDmrmInEDkKcd4SStDHxnlpPP80jecz
q7sytutHm8kN6qmk8V8tj8O3n1k37/ZhHAotOkPWr0eSOQepOnR5rph32gbUbmBnW6aIGt18jtUq
nLp2ip+lcB8lsW8NTot//xsA9mLVdLRdwYUUNroQGeCq2rXeyiELO1w44zrQk83O/dkicJMO5BZS
uE+RVPnpVN8QRxujiU3ni832WDPu01cLM6+ccJmuqK4Czw66gi+hts50H82b9BB2JPVsfgdfr+Vl
2CrSGSB18bF/eBE/O9F9dm4I5MqVb2ll0a1hx9I1X4ZVA8CQGaU4v2dKl/dt8Ozk6Kjz/BIK/8qD
ZwU8/0Cv+bbQuCu7pJFiqc0cQ/UgFdtTLxefDMf2+Dv2seMt5fADdPlthzrHFPzmuiCeDQft04n8
eEU54SAHbiewRU7O6pV+S0+rCiss7uO7YYZ5soPuOb8pN7Q+ddFAWp3FKLNYZXkAQejGnYWN/mJr
E/65Z06vF54MaOye5/vGMyV+7GUsdsmnnd4EZF/X1CKFcKnTddqcZk7ehJWVdWSeet9TE+f+AdGe
FFLZqvZzzv9+cFcqQsuTs5JIUjEOXF+/Yb6qAqT2CiEWqnVHmHg4SygTfo3DE/sGp6xTXOERXBNN
E9Tr586RIL/EnRWngT72g5isnun5VJ7/1t6Pjj+e2+8mYJDpVZlYojig2R+uexNUoRaOmlNTdGuG
A+xdSonWNUfC+niJ5yR3cZcahROlZbPurZneC8RTupSJJCvaa6amp0Lz8WnW0XapN5+W3Xw0PDjH
ToESLapnFJ88EQgVLalA/1c3qNZqwPz+O5ZWZMxo+IK9oobSljsE3zdHOD8q91ukuevuPT569kS3
GxdH4V58AsW0eGSVhKVDdy/dDOcvexYm0hPq3r2PYwghMpxX4j2xWVj16p4DRhRDtC7NBChTvyUf
ZyQuNpw6Sj9WOBTZ2X8ls9iIHiqzo+kb4FRmP1B0k7a57grwS6mqXIBTV5hF4lTQ1Bz0m0fbE1CC
DzxkJoYccRiUey73VzGwj9VvB2EUzibO9qPRag8br7jceBJG10nzuDta1yssDUNVhAddvl26eS+2
yZZktcCsLg6/NSQtrVYXiG6FH4ZNsbUN9slkVzc4fTjF1hDN+0SW98ta7wUATDE4T/YHKo8AwLnL
y6XgwEJP/de6ShihvyH+8/eo1NKljjIBEnLWBR1LU/aK1iLbqbUTQcIAB64VG7rdIGGvc3NFFJ4M
65qw6awnkR7Weali/AH1sWzz0tq6FJvgFIUILFYHH88xqGGBr+5Q6APJRbUx69bez7E8l1EWRH6F
PVqvbk3UQyyQqz5TrLv09OEK+pxOMZHrzBJdTRLv/YqSIkIm863R2nmcjTz4V0hbm2sQe2N+D8D7
mHdV/LIowsK5aldcfZhvDy5T6C9B6KA2uxlYACY7VQl1zqxtH3AJTDn0OsUsm2QL/xh9hR6bAwss
ius3Ca34oyhY6I9qshQqTk2WayFB+bgJRciNNrpA4vTGknPnNOFDjHzB7J3/+5+kNAXvERjlVecV
JBWg6Z4gKQiPS5CgJ41oV7tJYCTOvNVDtyD1m3wuGSeTxgyzX19YYYJAlpe0CTDuCJD2reLtB2vU
ojKNHoAGBc7TBULWpFO8v7Wt1Bn/jU1VijtL64F/HuG/GUIpfavBz9qlTbkNOqRea0jKDCmzPcLF
S20fhdno9ILGTyQ+hkPSkhDG7itOkvq/DSWgcno6bMaE2TL7W/f3OdKobYZJLAFKwL8JkqieCbAh
SQ8IfR6uEJgEfCwtoIdWe4+WoHZr/806Kvy3RZ0nTf5dcCNHpbrpUL5tWSSN5nPlUwSgZ51/AF5Z
QP8vlofzky5SP7g8paZbciCSEjtCzs/aB4hTF0NHQGG30Nz72XtPRt84Z5E3Yw1XUZBwk9OKSc1J
KC6RJYFwF+jt2SwEc9yvK1T0Hl+vBpbKUqtB3v3XmtbTWYhOqWoo0ZqFsCWhCBZCw7uDQKM3x8nr
X8bV/WtbZSZGolQjaiby1DwsPSK159rXaYI+4NSXy9GZvL1YDQq1VRk8DI/nRz/5IPIFa2DQAmfu
ceDq9DHJDGtW95c0B+n9BfS6aN0NuZSl58+fmxCxc7LXsboHpEnvkC3gdn8gYSYkxSEufLSCR0QM
4TrSBlmlA5nTd+M7LNliaBfSAQ+KBbKnHm5+r/bdKHn3zlfJpracDfxAUxV2RT0JjMz5HJh9R03O
9iKnsEOUHZJQm4iLg93xKbiE45u53gWYsb1LEOZ0Oq9O4SA9ooOeZZloi27aZRL9J4/oavi1tHX+
/G8TQO3RRR+y1e2da115moAsNGMj4M9jHdU3cnISvywTeca5HpvjVwVsFpL7OnMm0xzvQyG3NHiy
lUZKQVCn8SePNV71Q3Zm2n7D3TWtsCof0mOQP1oKEjADsFy5kgohKrJLPrvAsJharoNs9Wtpoy2M
ki5x3M49/g/1OaTwPe2ShJTtk9cwpd5E84SsK01UJNn5vt8VDu0w9KVS/qjCRIO3DtyAdZ2846CX
tdbMYNx9WGKXMRqgzbTc4Jgs5hVnATfTd3kDQXI94oc4k9K63XEAdvMiWzzW1XiLuOIBBfzFnRQ+
2ORpxA6kJLnoigp/629Szhe9fi1D6SOmUvQwr/VA3pBP1S2DEDTMsvI8KiIflgYZwTz3Ouf4GUAR
kFgSuJcPcszBcxA4sgDUA+s7nBFGqKmkdebNDRN5Sx7GBSZoFl8Jn4LODB8AozoZVstOgipta7ok
KxfxTYwF2BHdlrmwY6oN1lPASR0dAMSTVoO+bmyjJ++pQI9ATjtx1AfOZS3wqvPtjGtjx8zXF6S8
A+fkCxUlbExlB/3vQMdVUm7E4T5G7Zlopzw+plWYLLHNjx1qjE+XajYtZJ/lNUscLFVa0cKqPWvM
jOYiEMbnK8Fju4LnaTD9CF6rJQmRSXvNRVjbnZv/uiyGEMNHFzwF23H5CC7HmU6GyAGJeNU4xbnO
7AzYdWIVO8Os876CmY9naJzl1J5RnpJh7nS8LrM+smvy4lx4uGJYw+9VuFFJ7dyzJc0ZjMiVo/uq
oczlAqEZQAliMRrAlwB7ClibkpVW7W+u/kdpH2rYDCtDORIg6mnxqTeqwncaOSA2X70zdH5jSPBv
Ri0l8niTncMXMMcBDZv2tMRiOADUbE53f9LJQvsYEA+rCky6rIgfT1CS6H0kBd+5G6XFFTYRnS5d
tokPJGl4D5fzAsxL2V7cdJIjuXc1x8KIyq9Hwcb8Xk4xFXWWWEZfMn7vFEv137oiW0wNC1sySm3p
kYkW6koUbgSSv4H4utqaWheLgbgxUKI5eI7xcsCHyTYw3Ht9R3SK6Q03rQ4GsVFFZ/58NKAMaSVx
cXefU9gOqCABw6BGqyvJv5//SOAyMQnqdXpvgcrCfY5t5U9s/lt+VQgpf7VE4C6hCqkGB15/v55k
2J8chM3tATbh5fvZn7R47QoV+5PhITc8BGhWwPhw+sRzlChUuRmdLDlrUKqkbneUeHBwxci8J325
O4ua7F8+yV6Yok25yO+ltqEhQ8NVnZ8GiJW/SYJoDo7jqWtwYfN5rWhpPXm+UvzfYRvPTX7hWoKl
kxMGrAMTyK4QesnK2pZbJqzGkQ+Tri72UULSrBHH5VBZUZO/Nxzp7wiC8Eb/M5F962MhF3Gp7mha
6Lu5pVh3yZKugtyK9unx3R2W1w6JN48Hn0JYx1M2tSHuZzQU787zXXz7D8IbAIVBqq5/ragWx4Aa
SdX7w+00qEM00LAfJqgDE5PXs926PooBbkPjq/fOBJbqjiFv0I8/pNlXGavIN8PCQrnVAIpnanS6
0h3r3XliRZoAkfH227OYaiW+LcmzyBs8/ES/CGnTpyPRVheosdhzDSEGTiUgfDBjcrD5at6Vyes4
jHdlWhmzadAkyZ5r7uNxhOmNEgdGgTQKMHhthQXHqbIdu5EiyLjWWlmOlzav0Bx1DFGX18+Fu9m1
Bjhuv4s2veVZ4uiYRzpBSXx/rH/nJBPmQH1cCHnoEg0XxAOvocDu72arB6bPIwyym6HXGRPwaXpl
bZWOgqTi/Ev0u+MyQSAjZiGle9jJlElsQ55F+VpEsHXk9/70PPNzq2DvU4Iu52XaoO+TF4dqokVt
lWuzlF48b/0phDOUxDI1pcrRWEb5FDv3YLDjOTccxSmxHVXsiO+RP8EMbSJF1Qw0iWfTV4+BlBkS
quisvRWIWD8sQZ9ZRWPU0QuFZHmQcJNibu9S6ugSlDNMKHjMgdIZw0ChDYRExQtdSdIf5rPBHqam
YgzdDIOs+qGzTqdt79WHW4qneLAzn1lWNDxOfx4LLCnw3IhIJMvYVn2r9y18uOmOixF0dd7DpEFi
CYH3xjMA2GY09JHt2jgAPYUN6Yj2gTG9jllKnBSU5u65KFGsih3abJt4DSs12u9DEcdrTSfkovjk
1dgJgfdJRqgaRfxptJW5eEHVxoPB8TkdCsgnzdQV8S3x7pU0w7KWgk/th70B7RtIJUdIoQcwcnNO
QrVZch313cLKcV/4+2nODu0nI1Z54pmcQSHfU2PjNuX3SLgmqbkECoXIwxrcwa43bw+qGkAF+Kmj
+iAi+vzVMyxvRlLPmXA9wOBeBo5Gg6dVziQqXujNSvGmxU6R6ggR4nEfPfYTVzH28OKtbhQF4Dt/
f7rqt1l/FHxATa6+2YkMLvQN0+S2gA3DHZS8dmdkfH1Ll1BOvYo+kwOej7LQ5EMspcXlxV54/2hv
rnk7WISTDQIGBDFq8u65CbNOhxKEH8tGXRyc7M7qGUqDJkkL0cMNwJ5ZBuu2C9KqGGreu8ih9BWI
eIUIxtUb7iME11hpQMlu6IYYb0hAkQwXrPKuWN6GKg/nYv12bZg9R5enNs5q2lB4yBqbWtoSslbG
my0WV3/8cvMYIZccPR95beU+0liFe5dSYxW7IcxoQSvr2lQ7/IzuzoHx/4JDwMOyuX+tSTzFo27A
+JW/bW21dXV7wc1l8EgT3UHY9sy7Qv4W2PZldhcdHQuySnUq0ov+N7Mj+b1zxlT+Rv9qpjO360Yn
s8U5N+Wk28ODaTpPffLWE76WaK5IQ+RgvbAZXPA1+Cz289eO8e+mbv0YM0FV90hXjPKcw2/EYscp
snxl5qiAGTibZuYbaMav4xOdPbOAVwSBmDfeL6fsiCriHxrSKUwxmlKbjACrtmdn6iMWe42cLBv8
/8OpjlX2kAnEmPUd+9ufT6IeoXUvuQqq6ewK+qCL0h/QodYSHE0bOB810v0M1vDB6vegCOWI8r1M
wr4VR4TFWy9tAFUE8QBKl70U48QhEo5SzjHRKl2AUkQJqIot4Vkvt6K0pzt4btvCNQzEwHQSlVmT
YWBCNarPvU2K1ONZkySZp6C3PCnKYiuC/mulO0qwSb7wsxKPW1vSER078z0+onWUNxU/nOnp1lWN
otYBCdm9IB9EWbEylzInXVdZnATJI5rBoZ/JLgLqtQLyLc5mSOEbIzhLd0yaBCaUB5M0skFHOP2U
FiDps1lEH1wKLr+HA0Jwjhypuh8CsNsyipqRFVrCks2DFB6RBt7LO9IyT/NKpuqEIbXW2LwXgPxC
9BF2w/xUzYMGFzf2agNGSrYXTNX+2OoPhVoHMNHLqLK5K2QJqCO++miOyn9/yO3ZH+TjcfVc7Mgu
oZqpRDGLt5shBVoLm/ou5VjCmbkEuUVSRH1g7ulNDkxwv849L9WYdiTI65ykSlPVx4loS0fGDpaf
X28IuzYln1/7qELnYPbDvgpqMBHpL4/8GssmG853lfRbKpU3SGfL4Uk3lC9A1rDlSmqSC2NeYyeU
XeaML1srQKCMutVzY8i33ezvxFu89maV2CalGpNPZEMWgLp09XwreultllXpElExx7I94PAlihb6
WjR3x2EbCqDZVebkMlsXHryHYrn4CDeHrJivY9RClhXy34LbJPDln2BokugRoM6AOzW7czWGSfkD
8S3JFTyOctFc965SiVn5hwChF3snNh5YxiIWZqFiJCIGc8SqsNBpb53yWr2ekO61Y2mFx8K2b/rt
8D0pRQm4cea0nxBF/luNwmcgQqbHPoL7VuL29Cpyprgg6yUZ4mUics+w5+Eb0RCZ5z5TbS5Kzx2R
RUk420ttY7GAlvE4Ej4LMruN/f29TxyRtvCyQZ8ueQJok+zYSnDYUDIttsWDXCvrc6qLtN9Jaj8g
y72qcpQ8lDSVdeexm05lKkjPmlVCIKWYZz3HUBb/evk8oT2M7N8fwt0kvTM1A+eissk+UpKb4Z41
uMt4qbcWsy2k3GhI7wJM80BSubTrdjDxlKh4mjnlBsooZOsg5y7jFhkea9DPKD1AdgsBQ5c0i0Su
cKl1c3oWeMHqWVXMCvix9KFI4GGGRVeTO6LAgMu1TZBczst4ZEfClb9cZL6qKa/voZF1Meq4S+fq
crcCn/P6soxmhQJyBGRyoyfdu2JmTrIPci2wUbV1VFoM3JnbyozXDAySfUCX6pREhTSICIQlMtsi
mRrhs93EGlVGjrSg996e5T/X2GDt9i30Pa6rngLWBprTleUSmzNWAl8UR5wxOC5EmZ63zIwjdtYT
639cHSpMLdhI3lzqmDNnM5BGUwMmrKo4ODKP387irdvI0CirlEeXmtMf8s8Sx/8WzGsDvfIXGRD9
+Ls2QxRme2KVp+mFfVpw5teGdVw+1rj57Y2xgTw1ZT34tLkVJ4dr9mvRebh4t9zx55nK04NbkfAF
MOD9luXyqBaQWLJoZ1YhmRvzCyNG/ATaFuyRp9pHeS7fJL9BLpXfi8lLnCvhbGRo7pjQgsfT5WDV
0RklpZCxcmp669/4ik8e5mS14JBU00lF4r4dWGu/HyHHzg40QMTKj7brlyhY5Bz/bnOLXaUnGH9G
sOmxpYXvkvotKH2TpIOyCnZCdLQxYD2qet4dFPSyrHobfOJDJQK2YPmzl18N+ap7DXMTHVAI4YJI
1qIcPd+6KABUtl7tvCywfWEd3+4rLuzrV6oYsffW/1zXTwfsEQe4/yGO+HL28LhoiPGuEMgm7TPr
b96N3HZoaOY/jYUxF6Qfi5w8mi8/y10tQTpAz3OhD8v9TjRfQ2s9apMGvtQq9295CWgWnqCZFF0U
+gVdekprlFBw44E0m1NFDdWScjZB5F1KkGEw8k1SgUI0TLdZgJPZCaKuyqM3Qbr/ufnj9yyu1uz3
VjPh52G2pXXYzGWyg7iIw9Ul9WPByWXRoVIRAJ+C6fhCmtewxrcqUjPEvfu/V7mN2nb1NxRNIRg0
3jiuNDiRB5InBxGqnlMuSXvmsWyqO50qz7PLPhfE8rSFGS7inSOcVMNBBwuLHqj1R/7S9sFI6/JB
XTrPyNcnmsvylI8YygaB2e/kp+ZrPRSQ3iNJxTXs8cNlpHEQYpgzGOpimsnOXDfJ4ENGht8D651E
fc0myHrWf/p1nJNAvVTK5bDA1ieSnnmFaWRRDogzfVlfmZcMLr3B0DubBnQpcbLXPDdAmD7wlBzJ
hz8e7ixEwBd7dR/Knf216Q8aZVCm/9ES4+2bapBBzXaTN6pAiSKrDIctm0FjxeEdPtZCCULMluXm
twpaVstywItPDI+di62Z8LvAfvRdZFb+Cejet6p/NTJ0z7gaLyXTtlp4A3AyZBSGFHo6ue//qce2
oG1U6leW8x1d4mcCf5GmUjTYTUx5ls6ngTaHrJYPVctsZiCRU8Na9HoOjvvoKKK0eIWdn906mZ0J
Yv58idHdHpLDn14R86rftN0ZUOhg55EWmeqBBFp4sLmaduk4bVzIbNy+4Dw4Mk/WXhcBLMPYG/vs
pcIOWSe0S3c/cq+d7/x5Z/ukB8xmmMWNefOvqrc2UF9rPXD9kfXvfzmg173M6XNTaBHfPnjx2XF5
j+Epex2P6iGiQkJ4zrjmafB3qc2/Ot+70VdAvsYkgPfrGeWBHc5+x01NVkuRiyI6rKLErMJvDjq/
CvmiQHyv95HiTkZv0Fwq6zPXF/sSmU7BixumR2buMIbd9H0bbZnqe9kxA2gfcTC4F9ASg4bGvM/2
NpqhOuvnRt7lI5Cpg0hnM90ChR2eaJiU3DAqwAaVVhoix7gO38RsAS8OnoQiRoyXBIA6AIBCxVnd
RUIkfPmqaFLKcqhIquWt8m5vQKkqQ13mGQ3NEZ08+OEn9LVA0UDDHhDvhRkbnuOU3/j5bxsldlQu
R4rmcPihqk2816h+oEL7LR6D29M3Iu0OPteqIOrJZ7deFyeVK9EXxzWyi60WBXGRibrXmzWi4bpD
8IVElU4PpjnuLs0K9p/Z+XrvjZ5w4XiAurKIt/a60K9WP8xBQUDl2Xs587cvISQ0xkG4TETfxRc9
snqifDJwU3PDHdzxsDjwd6CSOvQHCoYtYzYW54NJL0IhQ1kp6W8pRP7aP6yuSh+xGouADPsPU1+4
5g6Vm4qG9R/yuMbNqTFEuRq78OSmIYPuO0yMeU3DbxCr5zX5FHKw1YeSoEL0qpKDKDumlWW6xvjT
pLg/1HXma+5DWUfwDcdEGtQT7A8IUjn9e+p6qNqJwKjASJlGauJ0gj6b+1IsBRmWNu9wAc3kL+/V
mFo+wLloQHCDgCACO+UqZGy+9ZXNGFpY2I/9c/W1OiJxTVRkldPkXM1F52af6vvhzT1nu4R4jxnj
mWlsbofQTFiCkIZU8VTl1VSl2RpftWGzP+D0gHSlOckft2r8j+aqIFs6KzNSYajgUQXBwdgsCI2N
dolQwnNTwPcemM+8HsnTnDY2hwCY2guT9mUPVxkZPExdSv5Esr6tHLMde8NIB0Gc70FuPjxFz5Ws
bGLe9D1wy2b/U3idaE+4HzM9xNT9jfW5/xhfAbVnV5OTT74LOIxwIK6xKyctAcAr1z6H2I09825j
ngy3HjsA+bsCQZygDLME+i6noYMNeQvbKfwu068tusWloN1ey0iJylAd6NfuwzvYndWaCHCy7y+w
OjnwqmewL+432WPEh0yrc/fYSlN/NJR1ATyoXm4SZihxGhnWCfT1waWyVakmP3c9/YLcRB1onBaB
XpwmDPBcIOG6onsJ0EIuvz55/BhU+COsF7J4qgQ/qBO+tUVDtuwypan342j0hC1F9OvI6DDD8Ta6
0SPadkub8RxsD9ya8LkCEezd2A3NqgfkaMwlVdr7lf1QjNnrKBd9czS9PRVvc5+sYI6Yaref7AaG
QrVBTByqEXLaVdLHdLSVlY2WWoX9lhXcs1yYiZIOBCuKRloP93X95GrimNjQd8+5t12l6a05OgM/
BsNaCU5QvP5aInoYQ3A2FpckOyJAs+EzF27KGMpUq1oXUK8/m3tJbq7TEY2+WzqRU6Ef7z/bVFUx
555d5Vkf5Bt0CR7nZduICghUk0cTWjseOk32C7k9AwATHSfZBFVJVi3crv9T4SNG8BO8rxAYicyb
8E8j46sN7Ob+UJlqrfwHu/aEgQFE1I9Y5MA+jpg/6wWwF5/seCx2jLRHSsfKvIXUTRdeZjdP82QK
a1V7K0L+mGluJ3iMo84nsgKw+SktldAxt7wQu9IUsZinMU7fWcE9Lkl5wIcGI5WxTpweTRnFkPxf
4Es46zHhUzSdadv3AeZlNCjlTPoKySZXT5Py2VNlTZRDAr7aWoRdWRnoHDz2vlno6iFHFpYSQZ8m
OB954VuzffCk6ytxykOEYn64KnxyTUhJEL3cQ5xv3lLXhhBquUCaHCQrIAnA/NJWHWxTMrdGDn6q
RVhNSPRAHVRqICSUimzUKhr32o3bHB2Vbl1p9fcAbvY+2aflQwvYvU+TZbwWZj1d0aJHhWEll62J
AImWzPMHFWFRl59fQXGksroVdOQN+oeZGWQp6t34r66vBl0ss9J9N6P4ucyPk+Y1PJy5/kH4cr+K
PBtKfba9MAd/dNL0KAWEKPmCN6a0Rz1QD7i2G6hZgnaCayVijBj3na8RW9qI5++NR9HZdKLCizfO
QsM2ym+vNtdvMeoI3+CKiE41PycrK4Rj8X/vE6tRJMXsmdCpfvZKeXkzi6E+Si4G23DWDleyLStz
eDBrm1JYIfHPW1jqKCz9xEyV10Sn36KSr2uZOimIGzhvFiU+UBbKvbCkvuFVkc/wQX+8UtzYX270
4up3E+K9gn1DSstbc/Dl7Lap76fXsxvJasgVh5us/t8zxS2/QwXtjl4SPUlaxclkvCq1PWpvRAco
odlqVYDUEUuLRR4gtEdFyl/zHZrWS2G6mDtEk9HLBZWFRuV3cewE4b7VvtHBOIPTRgCMzzkGcdoC
iZtnsOkG29Usucs9QeH3ni+cAMVZ5z46AdionnudDN3ZDp/1h+G7axIJ4aUQF1q5DS8KnKqMxHrd
bkytIqdQK64zhPDYBqAKPZ9RXbdG5l6+OXgkV4saEYwp5o4LkEyT9uImilIIdOCc61NNu8JG2pvk
aTDdCUmDJsHe675kBI+AQ8R4QtmWBxQrEIwtyH8/+4MnHq4BHhlnNk2Psz1ITra+5uFkmLUud/ZG
d8QsQ4kr2VBNSDYHXPgQmG4A4PpHZizfrgN9ad/ZDytkz173gRGVEbcbcpBECtcEg/hwlKbbvfla
XzVbF/Usrb+TAX5lGirFvAWNVWrivPntTztaHtAuYJ1hjxv1rxj9lp10oNz2hZEJIMj4eQWTs1B9
QEKVXaaeRheLW/DXINouZt1y/mPl7Y3PfsKW9lhdLl15JvgYwAvRUm1NLmj3s24SppY6nnD4JPTD
RPZQZDEY27au2TFgNLrYxMHugKiScGFRCokedsjfl2IAnu+1Opzpl/DHRjtVBR/CNaauenooKN3v
tavaEUhZ1MzTZjtOK9rD5XuM+/LbDw2fOxnPNRsL+RIydRyYSyOfjEKLvmZntBSHuKIP7IxmQyiD
Ce776KkfcEZAlAMS650k05wVLEM+0AhYs+6TX1TI/Zp3dqzaUuXVKpV6uoJPOphJ0Z6vsjBwjqfP
jgPK8Gp1QIroxY/OtXdJbG1RN4n7/GA7fmxRT2GqdsGFNZGvlKgGoudfgqNMLgrWKCuyr4uzhEhV
b3wJrp/dGeZnL+iokbZ8d0Nwj+sLr7WvlzshoJ92UyY9oAdbY/er5SBCG5d7BThB5BFvxz1/LjR1
YmIwRxKFIn3aiXiCsGhntYWb1bFGtEnMOOyh0TIgDvOkJudahcGudHGWjhz5AIFJkyU6OlY8MvQj
mQJn0vfAxLZqJ1oml1Qur53KWllEjVN4mc4KDFFfZ82HI6gsMomuVCvyveva7biDsCqsMvEuesIJ
Y0yOlQMSlEkb+eD6qCxnm0xMBqYczUSCN8eFt3V6N1u7MMV07UoSk5m1uEY3nN+C7Wr55hDhc/MS
gX0dbQU0BuZDVoWHMLaiWWcYj6QaWoulVlIC1nps4ks9ZMYPinYtQy8Z4CfEfR9SvceO0QlMwUp9
Jvb+9m8fNmrqrugUdAnKX2e322ShuzYvQ06GLMIjoLCul88vlIyVaXLmv5vYzKYIKsnYbILY77ag
av6H7/NCspw1Z4HLK9Mgb0ec4jh9zWWO/FpkOFYp3UGoMtxsg+Rwc5REst0u9PxlM2RrToe4Q3bw
021OKBeSTj1Ygz/UlSQm4d1+EMLvdkeZ9fDiHKQCW1uRVwQaw+KlDXvIGnBz3PMw1qN3OEqcQl0x
uMS3MDCYQSn+f73tNlweBFfbb+PQ+j9zwrd/AJvXIQCfCTf64zIC1yJcaU51C+5m/FNAsvBXVsBO
uIL4VLVMviWghHtx0LwyCWIRrRMcPyu0Q+h6XiiWZ3/0FR5xUBJ8CZDVJJ9KzlNaCop4BG+bJKBB
jyUlZiUU+S46lqCS6Z8jrGYbHaBrR69zny/+U3NHSJZ98cc93kPb88dY6NCVE1JIITdnoiz87NTh
zmSak4XAfuwT8vmeBJm40wo/yqIP7fJKI6+1mbrx4IPEKa/faYrHE3YLLrUWAFNoSXLu0A5tddkY
XqkKPrV6ZH088aYljL/Z61zK3FvE5wc9W53I7NfLdLErT7v2YJoSECf6U0GUStHTgLQk2KmYoTuo
5dfz4VeuU1L+pSadQ3IX7QSv/iL/aZSN3xe4OlGVcPG344VcaYJPYM5BK+KpNfI3WUi1GhfKXPxU
x0fU9nQrqpypRyunXgiSrxs8rPNwU9wOdx21PSbvrhO12Nh/sMWqu8Y5iQAxqQK1wPljxWZoFP7a
12WzqT607g4IaR3cbDqNWc+zYL6kgL9YB86Gyj624FrOJ3UStsywAfzpRbuZUPbp7l+cIiCjIG5/
BYKc7/wGifI8QudIMIVylJUxew1Hjy1wvz27GZ7Rmffd6svDn0hC1/tJ6JOfZ4Tdl0Y6gy7jvgUe
kNxUmuBhdc9tG/FzdaDnmRKPt/EHTZDBOP6VBri0D8KX2sXBr0AAzbm+zrrY3TJnPm4sCs+Nk/f7
vP/HizHnIb72vcYc9ZdaHS6M30OEtnjSHlEvvPIiCNlFUK34luU3fNW+Nho4MnUqHR0cWigKBWZt
8JMV6Vu5bgKfN0PLFg8DjMnnB3W3sKgHhiukiToVJYDu78uhKoZjaOUPGCdemFrw9ZBwz0A1Fr3J
FZSRJO3SlFvfKdmZWrbDpGL4f0BV9F9MJNgUFsHeOTUWFUvMwlB683fk8AHF2iVNCuwEKVCj9Cp5
TuxJjWE5Yc6Ih2F3/OhQt5g+ABBFdD0vQE5p0bkqDEGTCAbtWkd1+6dbkPgyJfSOpv5BHHTe9uTd
d2JmZoEaJXvTX7UgX3Cl2mzUwGVbaGbpIX1pmhEu8/oN6NZbrCzIAZFDqql1cuAy0yOEkI2n+Fxc
I/g65r7rXhTuNrQMi5LcYexw1EA4FyA5rnCioPGfSKzH6+dPKjeE6SDx/1yERg+GCz+AQ8rQP5ns
TWRntalDpcSAWXhcEXNZF+Y2n7sTFEm23UWjJytDdKXl00qw1E9C8/fJ/Q2B/koZCQ3CCVEjkLQd
kC/+h/54LyByAt5VKiFEEoWy/Fl+jI/70V9UgeOXMMogRJDNmwydHJKijcJVxThKTuA/T68y/jm/
J9hGWkX0CWX61Mhz9HUfH5/nPoh0awhBCNjzrDsXyD6i5UoV6Q/Hl3A0KV/mpdfUZgULoPTX0TR0
8k4r4uJO+csuNRwTCT2ulKjaNS2XYoz9H/+RuZl9mOVfJMDTbrCXysLoFqf5pIXM3LsDnLUSRF3m
pCSMjxJ3zBh2h1ii+iC8EeZysKZwT50Cf1FdM4torUlJoEUIEPpdyGmnVZWbH3C+F8QeLcbe5DQY
1VlJUyeWZNFz39mPBAtPQuu0lIMu3oufoXkoZEu8ARm2tvGmqMNHpdhc9jpPpgGVBnJNUqfIOHAW
uaqYZPfXMbg3JwGln3f3MB55rvmyMi6WrXpLEZZVySWhqOo8QHbsXmZka7DdL0k9Lxt/s9PaQu2m
WyeJusaGzaxRW/6pRJ7KpDVVVUEQx4KWba2a37uQ8Yq5Hc6NHSeHj2H8QxuSA9v8YWSyIgu7xHWS
0DiPMvqewlYbpOQAcBKzS80gbnZyq1UoZaz2dzh0raGyLWappuSEsrt4s+reU4NHTqTgluJT54lf
Wk+EL5I/khJohZA2tDjx3R2y6RdxEAB9NcR7Bwelb6Xt+X1v47icK6kfHA61WpckESlL4xtj7+r8
pPnAYrR5E1JPsEI6PZp3s3CoGmh1z+azj7CzQLdjVVES3DWD8eomtRRA3triuyM3i+l95nDxw+Gj
SMiv4vYGFT4BwXErYPLhNV11sGirZCQt+R+ICzppKSDyn60Bkmhk66+4ylNc9yxjocVuCRb6iZIA
O7xWGmN7cklFVXg8joKFDBoN2QlJPPzmNbPmAEQNOXdVk9EaluaVhwz5EFdl4REszNik12ymRGa4
sDt89zfup5vsWMaijN570F1xfXzxNKpgg9SkWjc3HlNkmzbb1yt7Fy1l42sflEtgpDhep82PX0sm
MdNMzCMGb/ihpe63HzDxKbyea/4r+XZkVCak0Ai7LyyUaK1wtfn5dYoGYOd/ZQ3qqDeUD0/1npea
rCXIYG3XDcccB0wI3A9PqCguOZ9FJ/tk0WB2IEh9d06Zv8J07WP3I/UJKvWRyLOInBIomP1EmzSV
iXBZ/GWYvdDA07SLgf/ppXzAP/5bD1BUKYcpChlmVrA1zXO+6BdaKyzjuvKh4dgNesIqFhgbOSXR
3fQB0noJplYTKHX/LtUtT1FN6w5tiPvxj9yNmPCIqrZzhshl/Hmg1PxccRqYkv/3aQ+1cGrK6thi
bpeEZCZrbfZTNKmNHzNnq/RgadkyJbemo67BXwJ4gSpRWCR8mMI878Ga+XBWAHAO1EerLUTbyCSx
wRhIj1YrqfTpeNPwFwabhecXHt5WLkcjtI8NFcdeN/ddScHlAty8fXM4o+7TglaXQr5eylfpAe5K
Rz+ZOUAJmKJIe4mjq3vUNBcdsfCH/vZ+aTxzOUknSXfvSJ34TSe/itb2HQgejWFa4qR4kseNLhsv
p2/92uK995VM3WODl2V4N7uGy6VmC0xRe40X72gAZZ0U3LazxK5wAN1CSqGWjvaHzXSZ7zP2Kbcz
bKb0E4gKNA/QB+IdxI6rzHL151VWNNJICsItazbGctw8iJoDrtsX92A7cjBYM917uGbNavP2UcNM
Mo6yJgkN8GeEmh7IEE78nRrATpn5klv9v+oOsn/w7VndSoIawxm5XKLOS96NriByCNs1bTmBGjJi
+7YPL3a6dZKcbcqQEV+Y0cgFhA9p8uMY3KzQuquYAj42Zw3ezFqGGOkTiMBm4w0HiAYIy7aOEUxK
pnTDnpYSVx2airkNJvgvOSWLNy6oB3lSMIFl6DMa7vt1LxhjS0PBk1mUpy4AyJUoAerxHGHPory1
jbS8Wn2306kq89d7449cwr4p1wPgyHX+/gB8GFrcIyxMdx0zrZxR+h3ZvmgC8wmSEpQgd7Vo8Prz
SjdDIuuc4y06up7jgykkSVOws2cTQz8WNmEoQcNsm6J34FXID2wy83+k2nA22fg+mHgMmr73CMVI
8muISSUzIKgc95OYnzsUCXJfrrkUM24lw59Iz9T1Af2CnczYNSZ8Xy8p+pwGIHEVNncZscAvSV8y
lQszG6JGIYwMdxrdX4juNkX90mDEoJCzDj4zABi9lH/2OdGNMvNJPpZ2Ikn6OkmM5ARxk/WMzb4i
4XUCFFShGcCFYzjKEAV1BAkIsLzMvmYCm0fvcw8TDLbDrHiEFSrKLCxt4hbmL7whXASfP4tJCbId
T+KNojGS7RXkDF1i+JnWpWzuzufYzDeOTTVJclfsNm/sPD6UUf/Hv4LhyyRSGq7gePzxQ1REFqqO
MBStRKxLi1+JjBXrHQt2m2Wybxs3wlZ/O3hqn6NKCfky+L81/Vc/qLIRXgBy09GiGqz5YW1Idrk+
BQ0w8ioic3WZlofrJyydcqPKzyQD366BWyPic8AtTkXHs2LtWaNCHMNc8nQiF87udxAortVxXNsl
vwXfa3A65qZcZHWhODR/uYklGE7XFUkG/bPJzASXHT0kKycYklzWsNOY8nCEtYurtm9o8hRKnDLY
VcncM3+3Z5H85rKLX9quYZscM0UOPqCG8Zq0TkW3WHr6r3iTDf3zauDWf/Q2uBXnVT0UABRPp21f
8pmWCGr6cejxnVHZg0+RodkCZANHCePtQALdHc7Q87upr89vdjPLGrPN44mpIfbLYyu6GSCQUORf
kROSPxMnM0EUh4M1Cg8ERiUyecALSJwEZrijsT7N8pfwJNnLwE9r8U7qNYKHkTaZLyzmbxZG21Jw
kGeUo5vtK+AzJYmqamfJ/EkW+vp1xSJvmB4rdtuNX9vqNAKdU53ElzgyaNSt8AtxY8wM2kC722px
DOXBGrk2W37dNHe+aEdpDotsQuwyDLcKbyM6Z/8h7zkNm+n0+/hONZ/4Y42qVL62Q2q9ruF+6RrC
bN+9mD8RhmTD1rWJbwzqqLxTbracPfxhQDGDErqAt9nK2yBJkDexfyaU4kt8cVoz8+sAs0+tozr3
tTpkO6Z8flX8vF5ftliti+/WZv3WUNEBu0dKmAEyyTqIo643TCGTd9ZDz49VZ4iFglXKwONuZiaF
nWybojXjQhzbLSw0JHuHb+BDyt4Wl7Af19U80VJ7bcQTWZ5UdiadkMDNqE1/Zbdc0Ln7fQ+D411l
6Fo5Hozjk5JDJBX2Xs8gR9j8hikqd4rSvl8X2qgrvolYiREEntqkWhn/qrPkME+tFZkrYAeu0gw+
L5oIwkSm2hVBY7D7wG3VFrqRh8VaTsqeu71nXSJEDOxdRckLjPhTaW5tNZUPwHoGsFl6bMEvxqtf
6EW10bgwiaHlsZsioHBrEkl9Iy+KZx+IXK0HRkZWT0KteV+b+R7vW7vxLrfujDi4ndFWPQifm1jk
GDfFmBNkwwclDyIP5uU7DCVHeG0az9r0EIWopJ8glzHYNT0U2Nk3LAgaC0bAx9AhSBFmD2XXfu6O
1ONJcexGtHgRuG1wThvVgdzeGrBfUjLMfnpv5EXD71WRgXguO37SMDiTvtA8esa2fpe2AmZxX6eE
+w5Qt49J4VreKvvCcfzfRS0qrDM7Irx9d/6/XO/O2itSJrMjf+YONpI1Xkn/4wkDx7BI2XGaXnNo
m/yGdC6iOvqqvDtQbc9F/xEhHwFXNTXIKCBraQcLoxbQLn2lunXerGptTLF/TaHHqqBQRKfFItvE
ud8mAxLFVzRaw9ZnD9wtBRyAsszWdJBwMHebOJtYoirWxp8Ga/8EqbTUYMKUFRuKUZtozd6G9/Ob
MDKjZq1LgraSse4pYSQkjFkQ/MFVazUXas2KiZNfVHclkEEzrzp5B4eevPVlEbP2KT98S4c0UDIf
Vzm3is3MH9W4DGg+9yT96t6e/HekBBELdBzHkJviJWMCqH0kT+O+39rR5FQS4Y3M6L4g5g1EoQS8
qax6wAb0trCfOLVKPldG8Y/EutrCVV6oesxqV7s/B6tysqWsrFNoJwaazwp9XayzOLueI/tbsw/S
/wSF7ww/8PjuN3ft0iCo1D/cqYqRI8exG9f54OV+dEgw9esXSH0jK2s8pnXdJcl+WRRRLJRf0WOi
X7EukxlxobmPuY880YKbxPdGycQ34j/pEtP53epjy1jIKjh9IZyx4E2RHLFXt8p8cM1tLJD0u7xu
n0W8+0wHYbGQZqSZAmv1RESHoqKSsr/jBNnQScAv/6cMtAVFF7u2QWME9G0suRBpbL5cXKbNKSqL
SjKc1jT2BCYTQSt1vd6fI2xEHpLiKUgEFC0unwpCfellee//vB0kF3VSUydxd0wh7fu762etlg5g
4fTZQN1LTJOyXGsnhHLEZ/BVU4rB9XdDiF+bVFf0yT/LjHoTOZg0HktIzHa4dhBIuQ/v4W+09zwC
poZXED8GFM5Y05Q0blhAizWlXmd5RBRdnnPPrwxKRC0Wu9bYoNroqPuDQH1LiBZYe1lz6xX0jMGC
fEz0/w+OzpIxv4cs+KADb2wqn4DGJNLtQarr6Vs0X3FcGUfpKhdaqgbCH2kCduahLv9CxcViDMyA
cgnXku5F4jmCKOFqBkLCIho8j978qblSGbx1QeqzDqfiox1i+Qc621qzXLoHXqoIXE0KTf20hD2d
7SvOVBXGDr985VZWeBNIkQ+hLjgDpDjTEQfNw4hrOxygMMoEG4P8oDE9BnOP4+IquuP7AKHYPQeF
2UGPf45vs5sfOuGGnPr52tlO+0wWPwsPkwA5O0hRhyCcmWteZn+/AKMqYwdsSs3SDOfo+LxpZrEm
JqFKgn/f+5T2Zy8FUhQRy0SpSu1oR0MyMsfkJCT45S1NsYGv3eIN+EIa4pjjQFJhg6wKFg5nupUW
G9dTjsehOD4HXdp697OELRI0B5Z+d9W7DOEkcgrYUf3OG3SFEEoC7lbbIVwUWQd7+XJz+QbcRE3b
QM996VQpyeUqmNIJfUxDcyj4CCZLHLozdD0RXvV1GvS7DRtPyGrcJSSFThwEnpfgEd17U3t+nafl
WzlqVhce9m+nzY08Q2ODkHcZ1wtDMojYyeKHDET7ZF34ImAdR6prQ8smwxR8HZjUMHTCzaT0jXUp
Okv5pd3JCxf2mcT5Xl6GUebFqa+9bGs+hk/aH2XrWr1wUgF1sFjXMI+j/OLu7Kvx8HVJWKpYEhO+
VS31rMnek3ZZGUdr9dJQNYvNNB4uuyaWtmtZE/aNc7NXD+sHgerlhBk1gVEI2TC50yLMW3XGGkCv
4OdFOocMIbPkfoIlwO30w7flid1KQXyWcAVJvcOS4CHLYBIJpAA00dlC/SzWB1iV01sdEZxi3grb
ADTrzJdHiUMPbR43AXcC06bAZ1nPrdAb+tS6bt3xS8tSmaA0xjp4YTf9c5N6yr/EADvxSsnwrL5s
Mn8PIhGHZMUdHzJvMV0MN6kFeBuP3wyz53xn7cvEQakrkdFsNpvbllqk77t4kUJR06a8jS0uULnd
cHIYXUbxeK/C978r92p5fvjX6Xw9Z3XFwQqph/j9Ah2oWau52A6DSBzM8yvirz7x0tHEZgU2qyuW
P+fRZGcFomjOI95xqxANxpSvIhdtSQgFa5+VUCKDJP2s9SGCoXSDY0/dGw4lM7mDrPwmcvt76dDY
XAhC/5DlDUe0hl2K4Z9PPNJztWIe9gcDAcrHS6R+/MqGmBRcMxU4tnhbJsLo4ge7/kktdOAUHN5U
0yrbH6FMCOwSr1dUyWHMnPBiUU2gGWYjqy4FCmROJ4Vc5me7VdQzRWMURZvjTPgIVVwWkv6vQEX6
9QZq5pA4rARtgSSKKLZJxvcK8M06brypXEot2HodhAP8rKxJtkPL9+U3NNGGV35maVDGBQIIIBGc
JZPkxTVguLSLF398UzdewI9O5E7J3zMUZHVIbf8hGVWuOwcsbaEJ7cAV3CN3f0SFuZAcea3NDMXn
Z8Y/WgOAPay12zG8wELzCL8sawyrvekE24FJEYpal1ofWZGyNgeJalQ59r9J/D8DT7mrK3WwDPp3
6amiqgsF+RAPN+zsp6JbqBpiNbzsonYvIOhJdy1tc3q11kYni5KE0+vGGIkVbj9d1V2xg7wHGTNe
4XBSf/HfLaKgbkqE4M21rXK50cvPAZ5jCfzyrjuTN4p6NSfefimaFaUoUrtW0ZkLObIaMY3GtHlg
4Ec0MC5Z8/Jxh/q2gsC9l9SU6TaCcyoP5Pl59hMFCX6HrVNbl1zgqe03MxzAjvYF0NUmWcjtRNTp
6L6fElqK4QwHSxkoGrn6bvhsyZq5vwm+2hP4aqfM7Yn/2IdYN/Hu7f4KQPl591R8HRYZO+lwVjb5
efRa+bzP/sOaIAkrTAhuwi47irxGsSS3+zXAW+Fj92Jbi4ZBCl5UU6ywf5FPWqEUftupv9rP9oX1
VTqM9xacymWrQBTR0EuZ5gY2wHSrS6rzpE1RR65gB8/O2kz+Heq4kFXW3ttL6xk6z5KdQiYPwfre
3nobGcew9a7tDwnrYEx/wodyeD2HV6Q6LED8rt1UJte7RGC86+lk2VMIl3MIVK6ZH8sqi0OnyIDw
gTuglMetOwkPdpqgC52RwrOm9GvvHKfiCRvMwq49qMJWi5w4FytmxNaQkVjnwIbOgq6NB083wEBx
y5V57Yvcs5N2sL0eLqpqxoVhV++JPOoSuDAc9RBwS1Ci784bNFHB6HVkOGSV6Wy7MmEXsQOPvLvp
fUPzQAAymOHwg8x1XWMRCxrpYATSCGGuBsszhUZj8sE2fkFL1Lqstw8NUOCXMuJHJiQfgyiCgB5q
WDdD87RfnNJGZFQzFlWVOhjaGZ2mOq16NxUvXO4YVu5m5KELC4aSHJ9FC2iQSXiBOpxrVDui7UB1
sl8YZrqT11+KqNpm207w0ZO/cJYRek1ls8wyJbZUzcknGcPs2/u3ONAtDgUqRmGknX2J0qPUR37e
RxDdrmeQ2yXQIARIfrhk+B82R7h4WqxdEeli2qDxrqtagtqeJqbcvWn8+wtE9Cm1sKwksJdlPptF
QHmHe+wWCKSFIDL/cPCt31d9SaH4Rkl1U7DW106BtPq+VCx7/RIhztZpieDSWvHT4+njYg/7/b1d
UnpmOAM8Hl2OGjYhhvLoEReitAeRAOHk/Dx/zJ3jJkuPsSc0oSRZOBH28GGW43OQE/rF43KbzdXX
ESRqDUUN8YT/yLtj1bXh6WCinz7ecp5cEyjyqEKt8klTYgv4cVdfXI5JwQaYoMVRBlFi+o+hBP21
T1kpT05sXqlsCwrdy3Ca6QuUqQLjThjBh+5Ix8er++eLBRdFqewRz5Qb64B7kT2hE7npWn+iJuf8
BvDO78tjfCfLEhFurhSHVwYRq1ucuainlEkwwPl80OTtcy1WYdpOF0qtPEcwpVQ/XB558lBdplhk
9F8PsYTEm6pcrDXyKdvTefs4DpjnBvwtaWCQkaYWD1d1pi4ZGPx5WugN7i+Fo8i4aR7680ZuH8ET
u4KhIjrDEuJCGLZXZCJbuw7SjDF5KY1hDYyKmM3CF8zj+ytO5Dn2GWiPWR1cXV28BMv1aqVuIUcd
GzT66V38ABoJiRwUW6RvEse0kd0uDi7ibbKckkTR4nuDcdppszSg4IUa9VqRtbMFZtBDnZuFAAFT
eps8VgZxtdP1zVbTm1+hri2VuK0paYIBEm5d52Cz6YMuxLQRQImHCz5p/dAVObKlySQI5dGYAD4C
bdC6h2WN+O1a0jReGmTUSQgKZ0Dfh8yC4sE/feJwvaez7JMJy02B717svzl8UoNoTAcZbdd5P2yJ
O0kZfwfz2VbYdJybjjqMUqIBwszBiflI0YQumJRieObtI7qDqO7DY2H4AJo7GPXVZxtF4/DFpol4
mF4JDse2GoCEoYFvrkKGy8cuz3pkNjh5hp691wHfRWKXEz0WlMqz8cQD4rhFdvNun5+wVlCM4tFk
98yoIjK/DwPQzWGJaAlvtjJXqrwuhkjKwLKH2tWDtQIwGFxR5vo7PI3i2d7La+uJrOub88WoYgAo
0Y+F7xrzQZPJ/uY9hC9z0FL6PqvMOZDejSuJKlDdifvlDwatIt6w55jiDlv+TTbqrqLO2C3jK7uz
fZejKePFlTppS4mqkuSqRR7lMdCh19nSzfbHKDeQdk3LkxE4bA3KLpDeQIMPVTodEJbttLfNTg8v
6fdtcHXxJ4CbjR04cirV4xo7zXhPSuL/nOR1UB4CY1q3pJKmdp0FS0bjphm354WmoQWHVPDVKD6K
l0as73r6k+qZ1V+tpN5CL7RjSaKnTm3p0V+UJaLA/cbPGPUJhPzJg+EBcW9x09JJfhv206XFoTfn
iSsgDPZZDfZQ9FnsUWxzExRoxnvX6tS6yY4XWvbtrc25+qQF26L1TH0SBuiLjv2IT2lB2DKptpx7
nQWOWT2jv5n5hxSlEE8rYv6yrd3Df8Q4hH/bXhGGMm93CghOxEvE7nj2Ej4A02PXT/tkM6I5hOxK
+HR9hTgagGqXAqOF4ywQKg5quankXnp68BoNhMHK+1hqV1/k35ak6uQ5EJu5izxC1EmahoOY3aK4
1PP/z+rmT8oQ+7io4lHyATQnUNTbDLr81pXGg34Zh+xaVkHa5V9oG8MkWE/xSCLtWQlKmOggmcrY
JuxOLEd//DlzrK2peS27knRtl6fE6l024PZvSnWfzmnRtE9O6G+0EZZVEzDqDxtxyu/ISfY0M5SZ
r1GukM6ZtF2kxJvDMxpDdA6oxLh1L+u42wEEnUx4qqQ+MCclwd8hgTFjomHZmyjlq1wYToJxddYh
AyeeeSRzpNURoWhIom+mVaNjsonzdO2OHl9Crh4yfyPS8Y4D3dAcpzX26CXi5uihwGtEvwFdBCH4
4QtKVBfVlZ4K0VZL6d/FY3CYrk+Ps/Kmgyntr2GV8p6gAq00H0B9yL0+EQ4qy+lSJBYlxOkJj+Kb
IkNAYTd7KzORfYTL6INd+fOmOL8opinZgN2YyCYMN+dsLQtgcOP9cUuJJScyFNnIgTkLHqpg/Eey
DzF9Fob3JoTyTvcE8LtT9iptNBziChU9aVWiDQpdyyUjS8bQfoiPN+gEZhoGNEFpxvwgC6+F9s46
bBKfe5hjcRYutYAgG6fvJw7XI/MBulwmOp8Wu8vLBP5RtN9xSyrAzIj1IdRPUfXHnypV25AC+c4e
kAty7rtBrFH8XCDL3+zjpQipQLLCPv3jPMzXnJsXVjbchxNsIRNVTCCqSyY9s2Ibsk2EB2x+/Cp8
YfjSytXzSguKKWDGoHOkQYmHRUb8WpxIFsi+tk++uYHd5/dJLuRsYBGrEUWTIRKHpyglbxQaeOvo
2oJn3r/OH5P1mCzi65BmzFg0+Y8T9T4j4yjxJ3WgxTg2qmyh7DWrHYEbheys90SS64zPZLz18oUf
SN21Kz21qCU4pj3jjM9BDj6yCvUyM29TFwNfGmvJJ+Mu2WGdft8x3mHjQDR14c+MWW6YnOQHrPj5
qaLozOBbbAjPix1pT5vR7x9j+edj1U/XaVqGqJSyt2ME+RigY1crkCql/OiH/c67ik1CdbEz1vbL
d6fxGaHPC5Ow7hFKlipO67KcvTkpXHOTXHniFXifc8KmmSmDltGF+gwpX3C4SMMhoCeUQ8sURCbt
v+87bD4+8NqP5LYAlnl878ldqJx12RPjYJrDFyeHyge+dlv8/v+K009AXZEea5pSrQjzTbwv81ar
KJ2xr8EMUIIz/jXtqTsuzCobG/DktgSB0ZeFOtdeMUO6sKa++n4sJqeh9WXQ+8rzuHC9Gog0zcDn
/WoUEVlHq2aJvsvhM1aiadbdd4EynHmJ8xk8onwcU+X8PlbL+dnyOFy+KVI38klUF17upjoTQVse
m6nvQYYMPwq+w1Vu46vbfm4eeCvOdf6wQlCsyY+nb2mOqVWbKBrA07+XaWwteEPBPWix7qEs6dqi
Lw8ReZ/hCHfCL09b25MOwDsKuvHzQ9zU9SiTItGgX1CnysZjCaVuM9Oakg3FSffxLaKgUwNnp0rm
LaiiaiP/0sbyQDF3Y5lOfGqASSEM7dvCyO3qANBikE9jYdOW0p6EqBBC5V3e+1LTFjCEObsH1pXE
Yg4J7m+CnehRQh1YypMptN0CA4PlZbPZbBQ3FyubR/XFotjReeHIbrovetM9VZW+qB3CFLVjxp85
B9ATohSUBl2Z+eeWqh5pS52j0mKKF7zoMsuKXdWoOq9w6fy/a3eXuooFnZijtaY9DaNDkMEd02Oe
7ALJxWsJuVMvzS/Qdtz+bsg/vwG1Gc2dxwJJMC3Qw7pt7dFlCjCouhotkV8IqXRluZpXMKHSMykk
KVbOoyx2wbH/5E4zvs3tmU4WzuzlXx8sQ7so6BGXo7/uNKgW6/7I4Udq3/1rX8kyIbooJyNA18vm
A7M3YxN81uaY7OlsI5AJR3SE9gSSqOw6RyUkod7h+qXI+FrxKb+JOavMktLWlz73qB+z40NU+Kpl
poHiFoHmpMH13RfpCYtPBC5usJckh+pW0S3NvYU98rzpoH2gBmeAq290tzATgJ6cHLDCEn2tgyZS
ZnHIBi2X50EXcWUlxdkimbI+BNfh8qo3WsDvcaUC9/f3zpaSesjAMWTC/3ktKwUJanq+ZSitt2GA
Bwg50oSCWjz5B1vc+xPfdaTWQb1OCSchLXpMPHhseSExntSfpeDIdlAU4PXiiOcHhffxeRtW7pOP
JrAlKE5yTXcd3FBLA8mYXI1Ff93EtGCy3AfqDt9qk72DORm6LTQ9Wpbh9kcEtFMfzidYO39SGHNj
qPSWLrtM3WMwOTeumIKci0vMoYV75d92SWLFrAcU+6uU84ysLVn22ipyRcPJoq767A2WCW5H8tdl
cciU0MYbxoB5YnhCu7qCYMxr927jCS2RyeR3bBrlxhObcfGVmFT0dJImUA0ZN1msaU755m0hwZiL
1HfzjMMPGiRZfEXuPu2mNshvSpHjmgJFDbrHb/CgJi49Qd/zgiY/jWM8E0bq/JC/fhSsHdnMBYCY
NJ1duKtliGjKRSXXXBtcPr6FlTxgKyyNiws+gw3vBdzat4DhJk74uDQIe8az5oN82rUVrF6VqAAX
YZmNadRieugcWauRYi02QSgbrply3w6VRFK1+y/9GWHVo69f6NQ87qqgn7CbaRtZDnxSCselpKqL
MzHDwG6Ne1l4qMHF4jUvuDB1M6YUffgDQlQpkwnTtrL3HrQiyXK5dYv96vKs1iyf1KKMl9E5aMXp
1oydOlujPgEOYLqzci79YTF34wa0IVEQkNdtt9iGHHbUswa1ouE3gT5Y3IZAT55SlGIn+APP0HvD
gymU87Bwz9QMRYvKQRf/HFn/+F2fY4YSOUtSQs4nE9y6mUfktEx0eIQrLIwUfS1StmFJid0DRqDG
7MSjjvHw8teIY2zrTC+p3IH/GGGRNfFvlmsZKn1ga7m+cDJXANBh2F7+yuWll1yeky5yWtXkPoyW
WbsD1fbfwNRcInQPbW1ZEH5/29RrTrYzHAThnMIeE5LASKxeiBxcbkSOR4IPZ8GwG1jPnPb2drGd
B/2jRFiKTmZWiKlewJOrtGVg7EuMOeO9McEcp9ngzcoGiWNonorpTIurzEg0a+aFKAyFQd6i3Jh0
z6xA0vuUXfdZpa557rcYr2X55tSOT3le0dBOiUocrfwWbRoYFFodNSLLKfFSrFoOXD1jNBzNbJGe
U3gdaw8nVo3a5hL5tpsCWMl3KzOSqiW6sciVRnBnyNFjxtVfcjtVLGWPuhM1ir4qn2KvBiEU/DSA
z3QuH7NRGk+0iApdiKoS9lsDavbPmeM7SlQCgUedMt0oNmXIk84mYu1mM6LBnZokuP1gqSq9y4Px
RAJHIDXF+ydAqjXZZ9xMjqYTm31nLO4qZD5kxGivCcv35JtXtmCNgH44QFRzrXkXGc99mlNiDAFn
PE1jEJ/7RrX3GOhOOAwQbHp61YWUTRx4zVBkc5ZeppEYdulckEp1Q/DjihBg+jDcp9Cv6w/sRkVF
QBPFWntbfCnuEcyfItpdgsrODc1D8xpjRnLFWb5uAq4Y8Qda+WooFNjMdc5Sk69wI+v7fMO9OOI1
qlXQBsfmHsr/hkxkVapEyqI6BxPpcYmWAAufwr2k07iddVpL92mN725MbcZzK/j8DDVDLoxrUtrI
lI3dO+s0jBoTOGzjK1vslOaTWLz+AC4DXSp+TAHkSGwmnUQeHB/A0JOaOe84Rhnrj8X1bVuy2AzQ
Fyv9xjwBZGB01UCtgXZYqVU4YJRi8BK7HcJHHksvxiERdQbVc6RnaGE5BRAR3a/CvMTJb13WRH8V
KzB8/IHWaPH9NUhWc1QyMY1f1PkkCXujhAneIE7HelBPDTT3/3gMSv46iesyuBIJcpfLXkS5ds90
Ayty45VdkzDhLPYHBfujwIuFrBvwZxzf8he0ep9tUYkgWya6xNeTUNfDOcB53Lnwlb7gX/+lj/gu
VD2WTXIJzURTmiKka70ZAW005mE2g3RYQyYCTQNhAExS80NGDRF8OROAVL6BiEN+VS5QvtvAXQjO
YwWvjJCGFIy4OUjGoATVQVZ4k7VTIRMvIz/uko3ZygUFKT3bDJy9qeFB2D82GkloU4sJSbdealIf
ZskW+V38LheFnlOlYMWNsHhKOacUxB7/QDjyI9U1CmbcqhGgjONBz950woE71uKYx1OzE+qa43Wt
WjGHaN8yUSPQ5ttQWA2VFw3q5ivK739Lvn4u8up9r8281Snh2MoxzCz6GZWi+wzKBvCKWPXhJprY
34f6ZCUGWUox/y9gB7hWAZSy7vC3oA5d8Q0xr/s8Ye/LvRZQ+qWSYLk3OdJ3mLd+kA+fFigdBUIN
iytfQJGDAlxTNgXLupXsncbp38J7Ql5VsRaACuUhzbezYF/jn+natHhL2lry4e4INCCEJOYQRJ2l
qmaGfP5yr9tR/P37YJ2c6FSdpJY9BMxe8IkhWVYS9iwwgtEGaSfoobYrE8NU9CaJVpCB7CXemA8s
9D9yDgMs1MkTT2yuGUzYGRgRviPYgGRpvtOaGI6iat+weSvcPrAO45q2imvKT3T+OZXSD52gU7jw
IOY1CFDJG/a3gEUwEgi8htcJklKefdUi7gUIaSyv62Tedags2DkOx5dVmXQNuHr7d319opEP5gO3
HJcphvjKA38iY0qkO0w/49jcZLNf/l+SOnv3u0Owc1V8ps1+pozU0v9+OlCqd2Fg6TofOeJpy9Xv
c6Wp6lR1CAECBhyWZ4KS/A/PtKfiDrxqeQdPaEpfcrj8ZSbC+iFcIaYUV3qjbfAnk0oQyFSU/sHC
3jqAEjA1ORUjlr9w1K62FqgfF0MnNwgCE8+Pm6+SbWNqs8JCvTWQ1+ukFpmuFitbap/lE7D1/+wz
4e3fyHHFWOmEcEUNg8jx7Mj/Jmpvlnkiw41hQVTU2TplREW7uFF3U1aJWypGbuUV5yJenxjNh+B1
SvONhg2/RmUOBMTmE1+wHr9R89ZPiOJleeYi2WaCtkeNWBWdFN7TKs9DnEruScdrWnbR5CPFS5Dy
IabbAbhiCpDvJYNl7xVSv37FEfOxJUClXYkW7FEQRMD00mkQ6QPJ/jpB0ZCeLhV6IL662aUkDdrX
mnDowDl4oOqn2RROvpuI2DcVvz+rJ05Neft23/mCt/Ia8UxGpB/bYsDTZiXSYpVkaxJsuKQ2Pvv0
xoRN4D4c4s1IwMZbqLZdMThH+dn6tVLjITdXHI4kqFRxmAYUahf8cCqesYXc9Oe0mabuWRdj7YAr
Cc9uEWX3GeTk5xgZhWdkn6ioEGLpgqM1WDU/tPeyE2roTVc5O5hlURrz3uQvM+3IVf2UXIFPzjJv
Gu2VCUUXroskPcTrqX0JEipL1FYICe7lvO1Wiz+cGuV2OBfXzoaHn8WhVG/Dsu2P8Td0trS6gjzf
mdF/QyLPXVaKklA6QvFagpGMF1MY/7DxTlyXplUcFPvdBYv2TVcc7Hme9SvrxpZV2p1oGwH9AK5m
2KZUREK1zv+YRZY5pKebX4trnbJDOrVxd/DPL/kOkmnJ2vBOwxXscfQaQLnGXjrmXfRNSbMq37PI
YuAg31eX+gk1JSQ0HjjYUxwcyUnmhUxUy8HMsko53z4htkjjtD4miFlNQJUqDWGyGcA1hHv8vBWs
5Ue/y2vQpidG/v/0P4+rp4jjqbplQyHeqj9DMRdu6u2dwqXeBFBAcUf236+RzY5ZnX0up51G+5P1
bZtTAGXPM+zGV63740VtD0cKoHCOgpDp8l4UiCCHHz3Mkmu/AX99ffoe3sBem3ppbU2zHLWmnT79
rD+j8sOIAw9fAXS5fB3Xq/dixqE2y4xJW7aOtDOGY2bWMAaHdzjqPMOshf2yoL+/LMrVKlcJAxWM
yxStQZnj+s+9up5f878wHNfX+oskr9C8VDc9VvpLKs+RupMmm8TbfPRTRG4d7DdxNo/yIJph/D+B
/IBsaRAmV0jo6a6rsJNXYTYmSECCy/3I/l7u5++Oo57srXpAUdZJUEiLIzgkrioCDInt3JygMETa
pnaBpGCYzxPf2K8yP7GeNjOJ9nOtapQ+0wgkR/0gvht4QdLRKOHM/NFF3R2vSQqY9CPhkowV+MUu
NafUAouFAPLAyEqU4tGQcVQ/9ZzdY5ExJvB3gJcIxkg6bVZZKfvscjlEt671eL4onAb6qDt76lRy
xYfbsug+zruoVrBWE5V/Pwp/bzUNMK0znATakVH50dMmMfmpSpR90D6QSdphdLDG2VVFVbL3NHrl
B9Si9ylGx0ugkVY3ftDJb4hsSD8CicBbauVBJ5E+zlZecaN9RYwWmTkiaM/pppQ19HiW0MkpEp9H
ghV2qMZG5eEhazVjtycGB+eIPxP9qAeTC2X5H2oIhBaJy/FN0afLeAMuBqWBMALVyTCUzXadGBBK
NbIOCO1fquEI8ViTFa1M68Xo2krNxoFCxBe2Gbi9cdO4M3OfHqILTLXlmGsmL5RgZl6dT58q7fOn
evJmZuNH0QjzVOvMDLGvjHuHu4ntlNKLZJbkwTU5h37a0VTxs2/xpyYH3jIcXjcp+1vr0t69iEib
iGPUThoCqT2I0o/q2WFlruZaqVxVtZIVVNvNoZTsiGeKlf7bJB+avL+uQ/RIO7rKcVWwg2P7+rLC
wm0L9VC44WsGrRgA8AMCTCCKsCxQxzA0+E7cAhC8ditNAEBPWFRRinKJY8d1PI3DM/4KXEjlhgXc
CRKllphm+Wm0Y9cFjqQNIeljS+XOfk/KHHfHQ5TOdfxkqK7LJpV5UE97QCnWbJ4kz967Sz5zfm7P
Aq8Y6Zw4ZflBoEGuBDCw6eD1MY62z+7QGFzVF20UWhg/Znh7Ahp0BpowyYL/YrKo30m8HfjcvMGF
d8vKrHV7K4/ienNWoD7DrDG4skD3RQDq8fiX8pCoTBoVtOtbMMCzyutuvP1GVqHh37GOnDCQy/P5
ZnoJ2xgDl54iqoEIF3i6TDafBTAvOIDmnT2lDLTB8X/3ezW59m7/2VgMN5ybIPpaltYP2PIXqtJk
U+EZnln/aJbVscPAa5rOcqT+OIbl9bAtBV0sxgjXjA43hRmcPU7ntWLsAftxggW4+A4va/5+rht8
RgEfxxzL9IAJFOo2vpe+or846cKWEWuqqmQxKZMSuvFEGSVOL482PGaofV2J5x9KosNuobTQTokE
cchxCq2zzmDMDtyfxXw8Vo6vsHkd9XvmD8X93ROgAWJ3utxZHKVcHYsNVe6CraUWGj4uXQkbateo
1xxkrbB2dOyTWz+Y9YNKTY3iTL57O4FenZXjy64f23R/PiFgfKrT44VlCsPU5xBgGRJlboZ3ON8A
R5wgzz2kZYbY8U+FSPrN9+unv+whbk5kP9UmN9s3lSEA4lORK3hJydZcjqu9YOu6gONf4bTyj5/K
j6hmPjmGbQevTSusezPjBefqKhxKpj7wU4A2N2RTgb+Dm7NDflmigfhw9HmqPFOI7XnvEajVJq0J
/88E5vXLU/pMN1y82uo/MPwR1dOqAqKOMI93mueReJTAmzAEfT1BNQ9HiQNXtDmWBkgyaDyr4JaI
PsX0HDKUCnq9I1DeNBJBjVjPYQcMpIwpeepUKxxZUMzbXozlydlOUEZ6GjahlCmads1kr7QGLki/
cWLeFwBLef/Y55Wq/aqepRYP0/brEaN+BHgC+Y3nHZTxkMbmLoGaN3109zg6Glkj3EEp3WALdTaM
tiZfE+duaehdniOeYZ4VkaYiFb4UuZ6szqZPQpr3UsCFXWxdLUH28L30B7RIwKTyC7CyD0o+FPL3
yNDUJ3qyxlECh2SM4hOO1nGW/90p9lkHR8YRdV+ddmX5YYCt1TOwZ9LPhvZ32N876kQdZBcynRqk
AM650dDYRxOHwe4+nDWf5mx/IXhcpN7IvXAWvx2qDhhsIlnlZsXitHNYDwOT0dFroQr1l+gs84cu
9Ftyka78t4A8S6kziOoSQJTZSmtmym7lVngAaR5DEjW7cEVhuk1FigkEBMKPMKNp0oNiE2z/sRq8
9YB8myogZcQvRPwA31XKAlTDBdosHrKjT8JjTq/C31CCJso4D+jxOjCv4rSw/IZDAMwfNS1BL1i2
+Io+uH4ChXi7BZTsNHpXA4SrQUyuceYtR90uPV5Ez1Bva0OBwn7ZBJCteeVdiiC7IUG2RbCbAt7I
J4tF53GKu4l1w9j5+85W4QL3hFT50joHBKG/ujeQYehnbwx9vkOJ76obYvRGw2n2/Ege0b1PHGN9
BuddOHgOBWSqX5e8qsg+waGnSD8CElTdcHSdqiNfCZfDuH52zRggiHX/xOu/ghjZwUqxf/xzhnc0
WRXwWkkBGQaaKqJ0NR96OkNwar+XZsndAhEoGhLMjstvw5ILvvGCwLT1ee0jfhHYu4XwIhnMFKA1
HtyRSTn9buqM6/nQxLw5fEMfPUEY0Z6l7sWybb2H9hTZarIK+iEqFgW1zSpPPJCJU817pGxYi7dR
2BCOtZLrDNNZjZmDgeD3bwhq36yXRrLc4vlf/+BnZVw0eNWDGNBZ03G0AQyQLP6Zk8nmwT76HzOf
ljFHliRkWrjmAfOEoTIM5Y3ugMSEnNX+5dHv4IX0wvyT5xIIhy8szhWHhFaWT4nIZSuVWoZ5NZ+M
kUMTLKZvkQ/g2qfh5RXCz42ZJk4kdKYUNg4NllF/dl47tEZ6mq0GI7cRpSXnCnj/MVvtXkqqVZHO
9rkvI4g9UXK7qYy4S+30tvEZzDNhxtZhujWngJ75a+A33TsRKO38VzcwJSzxSKQzFsoxIuUEKXqm
3l1FEHUAz0xR2e1i09/AciXcPWZRPKNGqm85x8AYTwWxHzsybOz2z9xB50APpfY08eMtvcD57HXU
bklM6r54e/ZFGJE3nH1TOhFOQvjVa+rr03RCsEBk5Dzowsu1M8dpoRUCjZRKUmbpdB52t5PGfEex
JoM78+KQMjiCQjTiKBVGfsufZpM9wBnM0ppSeQPBiGzJWhXy1x0WEgyN4VKgXCnwIA//shuzpErc
tkRlItKOHEH8nzjPuUetAFEDfD6IVR/RpCtCvOuT7Zkbl4uuImV/+kaut8LTNuE8j3f22HZPn94H
nTZWL4WQVgg3I4qaBZS89yfcw9yWvT8BrIgf+ABVLXNqeltP/tfM3T+0wFSpVxCA1gZEfxzREbsL
uMoihL4m76NavY0xEQy8Nqpody2ujpdrlrsCDLf0UGnKyUlyrH0QOTcEwSTnuy2L/O45co7bfl6o
Y9ohcNV1VHo31J1ppTVg26VyN4MlGzVoBxTp4TrH3Woqb9wan+6ZcW7NApG8/dCN1IrCwruBXbIx
zkBGn1dH1coYJOTuYzACt3o4SFEY9S/magiIaKHOrSmtTEvmxgWloPUIXAW+CUZV4KwYoGtJxQtB
SD21ENM0GsVOL5VJteCsaCp+6is+N6kGcPHFm1cm8T2p4JKHPFMfBzfCnonTqASzKfRDA1Zq2zf7
Zzo5VttOZw7yLVOoygoSPxKDzgXWZ4jK3euUMex0PYzpEd8BonUcim6TtJVULp+dS/Y/Bl6sxxWd
KWs0s5tSxnnejMwFQJn94PlsD0EddqCRF5pkMt+hoW8cW0z9Z6ThtLVOotj+xSqurp5Yt/KaGZRC
2Njhki8bwe9JQgH93aX5jQMHXP9RVHURyWokZKrf3C+tqzGND4zlodCRyvbgsatAkDPQngH93UYT
ncwMPx4w8D5U7B1OUKbsEQkcPM/OauMSpOawO4+wExRFcclQgE9u/iUXWEqz4HjWa04aRTfdgDiu
jCIraOYvwURp9Kkjhw0Bze0i8BqOcrW/ZRCIVExIfvCcas+3z4MSI5hjNZeuYvHDnHlunfZkW1+s
SntgPBNY7JWoitSs7646jBUpgiCRNbJygKGQWWXngO1uaDsbBmhhEgL97bKuaBEUMG0rXU8BxP5G
7y9hVZ391zbxfmFUxu2T8JE9xSaDYB1nQq1hZvlScnUy0aNZ101GrLpRVNyfSvTwSTySzld5TuOP
e/kXZ0FKug20NdO9V/sl9E64mmloHVyKVWOSeZxKm+m7Yu4+Au4ytXYxr6WxmWo5hZiS/L/cq09D
IXLij6mpoEbetr/eI16UmXDKi82QooF8DXC2p1r16zGhmfFu/ZyK4wzXDhYF7LnmWD242EdKuucL
ANjQQ9tfNyCupojtoxDZF41Cr2z3a7YTs/KraiY78Kp8lAn16X6n8JD7aTwaKXRz8FlcjHC/rsQp
GW1ksIqhqPyxi7FuJACjLm28N7xmLiD87ciYFTxzqzTvV1Hwh/Lk/3Z3Vw2t91nky6CwZ7XUSr/1
pqXL8ob6LptpefiBFBUim7T0ZJS7vxbq7cHc0qPhPHTlpEVoD8t620dJWT/xTSXL3H8nmbiB61uH
Wi7eQbR/Xa9atXswc6VGtDoTHLAPwtHUEdm7pbmynwcJP4cgDsQhwselrkmbMjnZnyKdTQhePsiS
KgUGMVxUHoOPeZcBNsz1QBnUDS3+EA+70pgospw5miRIRpnOcOIL6Wt+bXYGnI/bAPwN/go4ztnC
Z8uc7nb5QEFif9/UVvMlpmAVm7spb63vaZnCTru+vo4HDJtZTRo+oA4+wYqpI0DFgq1uhylVMyUP
HuzSWQCBJqTy/cY4vojXd21nP9jqne2p1sPMa81jMK13yyDYHrLqO09hWka083SN6ESCXXufYj/C
JnSRLehWUoda9ytMZ7hWebMnlX23a6IEermoSMCdUR5hT8hGML2FIGk2YHh7z8n4RkfdORRgF+1r
e3+GbvGJqFzCxdcLRImAykyES/KaI7xA9fbxNS67Za5ZgDooQHgEl+DLQFIN92HE0XFWfL5D292S
CpX8tcLfMt6IFIfoS5FCqj/l37DymifbHWSTzVwU87FSk8EhzJEWjCmxy3NwlJrLqMvQfrBtpCG9
upCE8RttVkjGxwWoutoC4UIAEDTi+hFTV/8Yidy1zfs4m3Xc2hTZ3lwGiC8m6PakxO5tPbmthVDa
avKpePHxcO/RnLH0d+JhAQohxKgVePvBYp1N3UyW76fxg7IWuOW9GxYaaPDVVVfE3W2J6sGoM4Mv
unjBCK+oXz17owKKPXrCoditJfKCo9DTHafCdrsuEd1dKiwIqcUXnwm6bdfbzsdckQWs4InGMD79
bRbQML067Cxp8H71QWKEVTDEX72BopV0csHT9xA7Ile1jHGSmHgs9S+ttrW0JE12ShSu9V1ZSZWS
JGnX7YIN5PysBPO+SN10XG0jYj50DTWNgNlaaA/PYST/RviLjkKC60rExnyi5eoh9pUn51ezWgci
5ni1AQuxs3loRWFQrOhZv+ecbmy068JvaxHDfFGzZbUw65d4xvCyuT9OthHPSzC8s+AqscjI8wUh
M90SkHTFhKYYRrNQq7jsCV8m7OxApowypEdDYDjV+KXSRN7espmQpaQ26P61xVEb72VPCiBlLbNe
AtQaUNODVOAYchv//Ulh0OI8sUU0R3cN7Fn3kkOEjbEtzIWjnuc85Uh2e5HkU4+ChRPN/n+azRd5
AgU6ufqFO2p91Uyhs3XaUDZLf6x9AkFuf+4rhmH4kJPtdbfz7Xo88Gu+afYzTavbccvtB0WYL4d9
oIh5XOHpY+3AZ9etASVNurAfhIWzhwDO6l6qgGH48rIB7F82HWGS5yaa/W7xD5wCc3czjZ+f390w
oAQRl4vgxa6BVFfFHVnAS9N+x+2cSrZM7uEuxSOXI4oeLo+4SpFuDXH1JePZ5gipCum5LtuehKy1
P9etBYkllUe96Yf19/SsiQ83oTtWoA3/Xjltzpz9e3iKD3V3PdeBhbpCFgD2BowSddVw+TmfP0qH
Ax2ffc81miQaqmHxyZVPXf5BJq45THG3ymyz1j7D/xuEC0g5PdS0jr8yq96Dy50KlGP+25AATrrn
wLtxFzG9UiGg+AUOu+5B+fARvfuk+U/P/wNBn7HDMQQX1salCLSG9R60LN6YzWKB6FzDjL31euU/
8HJru+XgJ4jzaM5cTA6WAl5W3FhR3Uuaidxx5kiYaM5GWmu0niFvffqRWj0Wu7vxPKLQ5Y9K9st7
3GCUDKgIAk7OaaJdEQaMwXaIqv9Gsfw8B0nfgiCvt1CPfi69t89pmpx/mhS+aKMLdb9GVH3Yz17v
Ly3ath7wreKLiPPrjBEK0qVtdpdqNkZglMPlcXB83mEKcMrIy7GB663T19SKnbiHJnSsZN7or+e+
lCc7L3yf+1ZE4JXzQW/pCA0CPRqS3yufYJl5Ht4vaOJiqogAKJnlS3cOt+GnfP7RvvxCOQu7EUja
TvbcnyZEg6Eot41SXFOI6lL6vyJqr4UI46UZ8DuzOgaO5GJs5RHFTiWk8Akm2SAToTaCcjX4i0yZ
L1iec26fn3DKulI5/+LGUklWpo/qnHAFbXDtNS45IOYLbI5rvCaVunF3rlvUnyrqAvSmmrg2uNG6
yqAgxBGdj+n/z4lGFHwG3ak0lDzRowNJTOfeD6P4cqc/TtvlmPRX5DDPwh8IOb+4t6qbxsEHa5h1
mzoDIKUd1vt+4Crwng8DjDoD6C6NhYfxz84mk+UUeKXnBgPlk5ysXYFdcUTfFAW9cmlewercSZhS
xmT6E7XWnpOa4481TAaSPYc06qDN9DfQDL5l/M3YgEisRsAWOUxB+H1kXmUFBsU021Qgm8p/0J/1
MwmSbYp0cUyW5vIpcUZEcuF6UzSPbEZhm1PDHDQ+9t/j0woKLQiESQLt+5PaW5sbfbShKAjHEVAH
94noRis/srXKYY9XjuYV5Q9qkrGLJdm24KpkZ2iRSlaPMBTALyoeFiY800MO4gGaw/iy1OkNqsTi
Vom685Mb7aLDQkeO8km+VW5I5z3LSUV4b6iU1R31nCFzYdjaiyxRcOrCmzdY17XUwE3EWHsjlH0E
KGsOIA/tytqvbThhit2V992jiu91tb9wfkKUtyWh8Nd2CUczDB7MO09/NnGRTsQy8UW4cnd/G40S
dAFdRi4gdvxHCdd89RhJCIWVRTlkkh89HV7PYwnZGWVn7Cn6qKGZxmRqQzBhVy1pqeg7Umuk9fF+
51K7yOoBLnmjymo9IlkCo4358ragPpJMD+19c5d5RVst2cbZ4AYNmpA1b4sz6FHQRtpQth+YuuCb
L4tL0hcWTochIlUzR5HsGQOvBVzEx5aI/GmlyfpvDVkNPaaUkdqTL5Fy8usSIkzh4ugdiHIlq2iS
FcbUvzJmSVMrU/20oshLbkw301uw1tGVQzf/T3Xl5zxbfy7VRJz+RFGo08S+qQ7Q3LX+EeVolZXn
5NZrkLfr1GvMoR0+UwY96bNWHCtNoyPVZCmosANG/eWRVK9BYfHCdx3loxX3wiP7OrtKxqPBf7Hx
czoibPUGL61V/+X/PBrF6/+LItySaq6jaZ0RN9ehAsJyrAmn7DcVwlAQ/Z+/6+e+zwnGoosZqVrx
2mYid4gE285ZY3pKwRTk7mb7Etfck4klwZFvcisPO8UC86XB04Ywp/fs7NaBYLkYbdIHQLvenlNK
ybLm7VDMsx2IAkDgZLXTYL42jams6IZ9HG/yZjwlIaGpS9babvgMbuhBxH3sAbEJ2d9xy1bLZ07A
/OXeKBqzN7GuRxFn5IRxs0MARrq0+nCOswDDAJ+pHpw3y6U4vHYHT69A8LlF8gzkhEreH5dh+lsW
zAhDN2AD6XAO8hg9pq6lk2QsgyzC6Eo1f7fe/tyHq8PmSaIalFBGBesx4pS7jqvrlC0xO8WR9cpr
yB8DoQGXVPgMpFRknjIidUaCNMm1fAaqENFWg/J3g9i1DJCxIykuFRN+Aq+slclmfV1IY12Tvds2
EHpK+LQNNs7QJqVGQgqs0jTTPK3n1IrsIuoO5Wd9E4158qOPsw+AVXhZ/PJIdy77vNvlh8UbdjNL
ChRmEr9oCBFXI0TyEkYX31iBI1x25JFggLIFsZtc8aoI11KEh3/vRu7HjWYGMSwHCFx8LANkXl57
SJK/IujNsbL4BphYXe4ZG6n6M/w2FFS0X+qJYyL9o2zy035yTRnRxtQqbi1sZsmvHE3B9NDtRE0H
aOUv9m05tDGmVlXtqGITt/gY6cYnnbAWOmSNE9qktdfbekS9ESf14b6FabwmuNGGVZoTNVUUDEVu
9dAbdZNnI5D9C/iV/o+wH4uN19/HSIzWp2UnLpsLmlvqfcLdBsE3nrfS/p3UxtZaIK3gqAAB/OE0
K/NV9sFSsOFNddUjxNur50GfeQJdgBX+fTWoAxzacgntX5VyWOY1x6TVuUel0WIzUAYWvA+8xhQ1
10ZR5KpUxdZkNg4WVGRLzuV5rt+6CcgJ6OVtbzCdFNmH1avNKGfCsccFYB2sF4WtrjwRpW8wwQ71
oMHTe+pT+nAlwK+vQt714zsTSSYspsWXdCNu+p/5s0GUWRIDqlAjiSF8X6JNhEXTUfVnTJNod0d4
C1GCrcpgLTOQtaN08mwgffcb3qMn8SACQ/MnwqXAkGUzKfWf7ZqkiLc4CNNAG4iO43S1eZH6ep/r
Kab5Lzc6PP95yJ7DLTqi29eYgMYNZVlNOXbTIkowqk5hgJEjHvEGpSldTiEM+215GWjWLoR3R1sc
6tYBKgtQJZprTNjBTktwKUbeN+x7ppvJa0BjTRW53ISF08ov15/aqYdujPyWy/jdz/ZIHJSvchCB
q55VOuWwzL9G1UqRraFEBlm1nIWwAdWIaGmTT3x+SAZJYzW43yzcUR/Rn50swrqWDZS4Xyu7iPkc
hbAHjII9C7WJrpzrPsJIAC6IdAa3X8iJU8r27TXxrBRMsn0Y5/N4gJ5DgExCvKT7abhT1tkRA7H0
21HzYzsXDSMdCms1izn5WwvHxqSI7GWkS852Sbrs5p4dms6YW2+JcTLKc89DaMZWDzCAlcE5ud3y
VEj+4VGcoNhnKdxnjkJBfBEmHKPTfnxm/aXYTUi5ZlHh3vDDYBQZ4i5TBm6KijYVt1U7UNn24RXq
mmcHqx5/UIsR77GbCmmmSsq8JfKDI4tOqfNx8IJKeUtd9o7t1ak5JJPgSupe9l2It0YBfX6z6kDN
I+JxSXgO+4J7K2LmAhA1yL17nqvi3lGYTX2764P5CL8J6mhPBq8fiLMlY/kWsoZAyKJ0nU5XkWmd
M4cMC0IMvb1QSpCYQJebxJiFjeuBK39LG+IqDgf4gC77IqS0Fbm1ENDN2WDkKrgfQps3OSTgvWVz
TsD3IvUyK1j25wwc0MdPDVG6NHvqzHgeR5Fv3dXawPxZbslV80xYbQn4vL2BfiMgSZhdHLu9FeKU
6xjAoI6mS33Qhfa1xuv1sBEGz2q8UXsIGcJCJqQzC0+Sue1PTQFSDmqQe5LN0wgh0Y5xiRDw4EWl
EDUtq9tiMz5LvBc9suSOyDBtM5ingiQtCaoW6xqxS2ONHTIIq93LjmUzLiSGU3ZeaP271XksuIGJ
GxZVQ2jcpjQjtELn5o8qP8HNgUp1DdU1HwF4xWYyR0lyfoBRW5uMg/Rn3znCJnCrfu78y8hsKs2B
EW6SeZvaIbPJyi3PFBRUlQ4wHzN3Akr1UGAbxIw2wMtmR6piqm5m0IvMVgZhUn9G6LWW6bpOK/FN
9hEdmj1l3y2pDUZONHg3MQ1DpnmszltQFCDJElVCImAgm7UqgMPdnIKrPU75S3rqUGkZGpRahAbB
NYuGQYKTngo6Nsn+i4232dpb0XEdzl1Utsgox8sZLXSLYTfLIVSDmImljzYhs6Y4QvTXDKXywbDK
I4ODBnlmL5vArKA4aEUJMH54W2uanABvSQgbHuFi9/uiX0cfoTDV3g1anZ+ZkMZjZnNk+Xs/A0W0
au/Yc75SRDKiB70ekGJOgdCrk46Wczv1RsN5e16C4GE7li9pyzVuL7/ZY/qD9aQaDzEsOdS8+7ec
FjuXW96BDVaOiWLLQtPnZmrZ4L+sSBKTCCLlz+jvqg3+vp5YyPwbsbGjmS0kETiPaBA/lEjipytE
JzfqCdwRhJD4DWwy3CX+4N3STsFXKum+tjF+Is9MFIkEcMM37tZKPaN7feAZ8Y/UQwiRiaB8vNbm
1eokatqQyZ0gqiMTgESgDknE/5WLRpNRdbhe2C8AHXXI5ZPQA5SrI8eiG6HP3n51JdZ1SNOSyuW0
MwFdHQ2K+Rzz2teEL9agHsiI2jT3PUVbk6Gyf+WMDeSYZjUD12DfGQPMs/QzIDk2AtSe7gGyfp0q
jix+qWVqj3uIYgP53Epr4LoG35xPAEd/GhkqsWpAUOQsym6TRmHN5cSCthlES6eSmUmjnK+i1bv8
8cNrP8u8qxci3YknAFRZT2JZjnabShddZ076zuC7vUewHA45AF6G+8js58/Ja2mYgtyUqf8003oB
e8CKtiH4b6c1cnMpTmuxSa7QUdHJXEykFiuffu70lsCtY+PCXn5GiREo5b/6P++KvfCyxTl/wVk9
0HpDZmvqc8VUbhY+Ps6fQ0ugpSxGXyT+DDZmMBGGEAYAQiyt9eVosC1Z3BpROOmmwgUfanqjFjqz
Zir0AJeJ8hyJwLRCqaUYrEf/BuhcleTUYmbR+afIH9L4VBF7rckAL8J6wienYtnLjxpG6ZgHKiB3
WI3qmw0BZDpXkVFLlZS/RL2Cv4v9yENEHmIS5M7GF6KJPcfG+62xN4gjvWKjZ37M5+9eYYCrgJzO
PwBuo4Hw03Ij1KeBQSVWZXMyEw68rwqElsg11KB8bEc/GNxkhJnS39tSzllKUNdsY3lTsqp8MpvK
o9JT6ZM8/TdTHdtFFOw6PpVbM8VZ+SUcB9jSKTUr6hv6LSJx0dl7BrLipYUVouysgNuBn2xUYHE4
A1M2JLLi/CYnJFDavjtEQULLBrWwcEIS7Vo06f3aD/mUPYR+NtUA6p1NZEtlSBGT/5FrTbcIG3q7
0JOxwfkLEOkYiW5IUDnHv8tLNnBQrLDvkBBMTO+xqiUHSn5IaJzXYlL8/oFTiucHS1z8ZN27zlqv
soRerW38uIBfu51+EuMv/7qNUuUK7KqYUHhWYULk2hXK3xs14QIR/94C03Fz37QIzcHGPPDrAzzw
8DnRgzexwtW9yNSnXdRP045dGO+S/ObJdh43LT7JksyK/D+NQnWI9YniBt0etlzEbVRi7i9yigVR
/udjDR/jQi+solD65jscr/qnV82x14YO0Vd3dfJ/UWqz7sEmpp00hl+oUJnYXCk8OaKQ9NVupNHx
Z/dgQH6t3CTJt0Ymhub1pYKLo7uE6A6dRk/JYfWY5l0iVfKzGzTkfKpVMfbfxqzSE3S27jXMGREO
9N/iHjkLrHSVxqbt0sguS7Rb5M79LgEv6uvVy4aFnreluO20u/9XafxhtqHcRjoHimX8fJqQmO21
S//d2wcrf5BRmN65AfRy9hJIGFRy6f6E64aP/eraN67Hw5g+IQdfd5gCsZqi4Vf9tCeUxxrb+FN3
GRukYU0jvsjEJDK7WsDU4cK7cCTgP0FFqA8WURx1UlizXGj1tjddZCc1cnbCBkFbXL9o6gq+5dTG
teGOJ9muRMQEWpd1DZRl6G5zn9F9HHzppGLBsgExPOTHbIt8VIJbGWA1w68hfFgag08bdtxk+VpC
Q1oLeqt2txgg0dBj7za+dZMINKFhjKhqdNLB1W/Vopj9s8RR3/FzUdWooFIjR0q9a7nDbftlqThA
0qJHo/Clh+Bt1WPurfyRXap/ETWOfw2XVyazI05Dobi0HPxwuP8ZQWZIzoy+eTT2IesduYVlSZrE
RLYMscNsjf0WtUnLFGh26ZPwp0c8bZzjyPz49LSFLke4wviVj+A/RtElCPtQ3VsiugUgK4fXFWdt
fvr7TqAdHT2kIeIqSWoMcB0nZRMZYvVpD9wyGqqGJ6A05gtteRUBMAusiupRupwLUygAtMn/SufZ
jcKCO2N4PVW7Ktn6/gm/cFmVBdUWIteOsyx5Gx7YSqgdb3SB9iJ7JFCwIA/T8IRWTOyDe8zfaDCg
9RG71iMmw2HoMD98RczHPKYonrhrO4oNRE0ll1b/tEgYzOdCaKGoErBSBpwnXyw6UVHjpeuia3MN
dtbSjUbM91qACtvQVFcFcxTN+d5AoqyMbIuuEznxjEFs6ytdbb1dJeS3YfDOA0TOByu+UzTvx4qd
g/ajJEmDx5BgO/AdJbR8G9WuSEAV5ZhYtyzWzRIq5UlMusUsUI3dtHBkQXL7l6whFTlmT2y9Ekb7
5yyUhKdAMAug8NyvJVv7gzgHGdDZjAad3W5+DJqvfD/LSwEVs8C/VksdC+VecfuDFY1htFYm5n58
TiLd8qoJXDbiHAuzE+6jkMkw695Yn03F2LDN/5z+tRizwAcl9iDfNqvL2Sc0RXJ7KQ/gLEPUiiES
tsXRjZ/ouz7+wx+6w1+XZNzRQn0iw/E78jimUKmgd8cTW4iHO0r2kh39NNIBTTPl7iqici206BMb
okFyn8I8LPpUa9ESMv8JcAaEkuHOyzkjetQt+5K8ntm8tYdww6YOrDGUkbV67jR/aqdJBST01yx4
2++hGXvwHnmTqgvRmaWLP3YYxmnORmecX7Q8zGsonaVpNlGP3quxDwaM27YWjroBzXRXWUE9rYHy
BdY7lU8r3oY0L2fVUYCCFef0iPxqy4hmYhP+obxkTnOtjOui1O88HzD5Yv6uTcyG6PAs+TRNknrB
KOfkP7ty5tj3w992HfFWpPPJYeHPbV+oZe0sQlqn3NxoTq243I1CmwZGuPr9SwNaO8JKYt8NT3jF
/s9OtcKFx9kF5Y+YfVnh0e2aG2Ykhf9Iy2FnHGlqg5c58o0TK/HQY/E5MedllM3OMN/4pSLsy1R8
6D4M54yAZXT560BmOvYDSFFxt/G+CCe5L9td3XvNNpWxfwfTSZSUTQZh85xHWAFkCt5jCZwn/l/K
5h7Qf+FFdb3D+mwck0IcEYkRFxgk9NrrQLuXfVGACYfXhVQMeqVGjakDNpFlUZroMW3ftawNKx3n
wj6wyzSCp7krLtpK5T1ApXK9cxeVfodUUzq/UkC7We+LC/gMf+T3f8HBN6T7YxrqbY6hG3HgIZQ4
dQkAkUUWoFVSqT9qGxFdOw58VtSTBdszPhYkC1t4z79sIW5UggLjJbAddnXH3cAtDZyiaqCHboro
hXCQr7DbJv18Qk4owUkRp3CS9kDivJhMCP9DT6C7xp1DyNrvc5T2uzbY8Ovd2tIpgixlcmBBmwbY
01p/8oRyEehZ9iW0hSkPDSzMOVh3FTaeJxmJKJdWu0Mb4bKD4WGhvx/VAacnrPitmr8Tt+JumcLo
ueoA0iIrUwJavLyemDCM+KLkHFyffeeE9iVKAqa1tGJogHyYzg21E51V39VRlLyma1g+7RTR2CpA
bW2teJGUkn3hpTy2hBSNM/as6kXhrghv8i0waQWLlTrz0r9iCdFl21jiSQhw09EGNX3W7pXbS8fP
0hxF3QnC6agTPCFQsPB2o14HEw7kHO6wgzFGS44cw8onAgNgvFn9YsisMxsXQ+e+RaE2zuN7nnzS
Yk35jOpfonkmxCufVAi/tJEuywAC4aRwxxO79YgK9/TciCdmEVMElJCE7jiR3eZV1ovdV/xdJLAN
QIh/4VVD6szsrXjwk2BEXId87oIeayPUmfJtJopX0iLrOJZ3ygvAvo8QGIyWLR/hxK26hDY3SAhT
Xc8L/Gd2wQ9eXAMaeaqX8+6oQ3NWQwfy+knONDW9IbO1QWCU9QuXnTpeny94t5yy/qVl/ASc9nbN
+OU0Ly0IqrLfjc7kn3CCstZtO0p/riDeqm11QJY3b9f1ZYwbleBZb9kj6jC9NlFH7NTXb+4HhCTY
tbKECVoK32U8e3WD7oJA+jFf95MvuQv2F0OUxnaMpztdlNnwF3V8AJdstPcH/uizgRlsYQiDVTHZ
5FO7wKR3BOtwHB4TAGp/iSu7wmPQV42Lxo5gUPyDK89QOwoar7fYsRg5bmlDsU2yWmdgMGKm0XUn
zQVvctj/OAjU4GNbJM2yTDRoFfXkIojmV1kSzFWJvI3V0lURv7EaATmH64pmXtAri+DNtO8NyG/f
9Hz+nYBRV2Jd6zkJ8wtwzLZC1JpFpWlv+vtb+9jmlVIXSPjnE7nAqu43iJjRScZyveKpdBdqsSdg
mPNCd35r9Jz3id69xMM5Wt/9oJ/ak+HeXU3mGkS1FH1eGc1Agp1K8UBql9VOPgUeVGsps0lhfIa1
ZMlk0cg63/XIQBRnudeAbEtgQuZTr1Wdk3+bs7fFyOH60o/1w76wxXfnwe+yIv8t8JHMEnnh9vRB
qH5C0sN+8JZwsZex89WvZIdeKvasXAzd8lrEFoz1sYWOKILvX0Tkzeb2TX8JTMkzHAD5NF10wMNw
l9CG9u2wf4/X8w6L0NHtaTU/gDb+uwBBJOC/Z4WGocclDhCY4O3YeTYBEy2qo3oy1Aw2+ancWkHe
yOU7LcLglnHsv9H9OocNksl47SE//Qox0+PylJoL29H1XblXrQ2zcdSX+fqBM8gQMsnv9rdHlKtR
5ITlRPU/PfuBnr3b6OqLU9y304tdKR9M+OrehAolP1bIhSjQxXSCgrSSwWC+Ld2rRazR1rLH2B4u
eCjBP97+mq1ERYbj+hAcOD/fZwdKcEHSkK+XUPFeqUCvnYucQQSdgnYTjCypdp9/eBys8PYH2lMF
UOmPPIfLyGYkXejxEGbX0RaIRSlytViQlISs8GMMltsOQ0ldEVVgXE7206L5DNZOvPDxAqbu9MuY
K4pF9e0ohYSokZGOYcU1nrqeudnpHvsenplbEYAwkGj1+FXCVJ7LoFjjxWwNupQYT2SrDNWn/JzB
q5L6CxX5SYZLpelhaa9yS95tB1/+1+8LR0nw7miTnVpsE5FTIsF4Ze59fcLuJuLttUbhH0j5MtDs
jtYZGSXLQmdhw7FkckJXyi5Mt9GADIOJdnrFQyDQQKoHPkf8fTKBvtGcxRHBXjzV9pFinGGJcKao
WvQw1jUexHBLIEDaceZ/j2BiGq5vX4n930/PF8/ANhd8t8mVyg+kW4zjPW+wkY8wK9tPFEG1l8QV
lnsyPJd4iFl6K3st7DvMMZpwnAdszCjk7xTTcQ/y0yh0r0FHtexi2qCK7jrkCXsec/By+euVknN4
4edT1UIq2LVs6ndshnA7h2zDW8KYT/nfLP88QbBCWuL5B/UN0H5V9EnjCAwsPBmgo1fCymDABUdy
VKv2xCdkr+BtGFMMfaxqGcAU09AhRpmobHmje7goYL+RQaC5hdgkWoECaehZzHzlfevf1EPv5wlk
qOYLH2EoaT7+I1kbz/wMTmc80IDQwsJPLu7IFKGqrxxxsmpPmgjwy7/zWYKC1AbCYmxep9uMNm0/
5Fxk3PatP50dSvl/+Vn8AJsTBcUjGa9k5y45HUDT6kCAVngsaye88uwRQn/bbYvZfwmC+ViCreVh
lXYU7sbTkMwRK05NVa8LsGBfHj1KIolLYyet4+0DiAwmZ136MTgo6lj5NJ4YoaajKXbjy8q4By9d
NDM+FeYix1hk4f8CDcOfEIs9nmrkjypFD6QatC8fknv7tmIPsU8BNPg282lm5TJvAuCHaVrNquio
hAmM+P9cemWgAcVIibU8vzhhpI9Y5NKxE/uwpTBAXyd2mJ1rfYUtZMzQjLJX6nnXTeyeEKbVML8W
loyyCuyOjhpacnGVXIPcOVqqleezkbQZ0BTIliIPS8xr4bC+GYq/KxofGmrhjYh+GQdb1NxWk5Ih
diwT7Dqyr8fQNRz6rMNBv/sIpOBpiKDn3S7G+JbZxahwp9chkqifLuTGQbirroBY189QXcJ6th4q
r/bGL9Rwd+zr6nA1BkoAEuvXLyRv0NnKQ6QDfimqvF0PblHXP1g+fox3Xqi3nw9d4NJDdMhxfwIW
7ZkIxmIDZmRZ3s1HxRxDlj1P/dFSwbxdjTDtNe0QcjzWaVpIHG6AzxwsReHaxq6Hw66OVlwRgJEv
4Igh7LQjxCAIWtHx0wPsOAg1fd1mDJjRn9u2e+1Gzk5lpZFaFj9lrLjkHWcRu9ZC8nc14kud8Rby
wQSPzjiG+YhC2w1HQEbcQxiAS/Q4a26PzqDDkhHkrVU358cY0nSwBPvERjJMRTkK8kjUKjhpJWL7
Sm5m3LhWd+NGl6LosqRrr/EDyp/N4gAmo/nwIWnBeVwk7wrWOCIGbKzSOTiSdbBijIp/3hltega+
jvZS/CZhmadv3o+HyVOlxeMdKJKJuJobti8pRqbQWJyfgb4h/wM1owmOFnq50U+VdbI67mNe7afK
geYouHqvB8OCdoXDE+B67vQvKYQelRm/i4Qv9xyW4HVSIsm8G8s/jdDk0uq/KJXD+e7bUVFb8kpR
HaE99gUliUZlImN6lWM2MK/2jd8TWaf04iL1n18hZJkYNmMS6zi1ZmVwAZBFOKT8O2xH4g/ChbiE
2lxl8yoBeLYgunY7LeQX5acP5c6174RDjTXLuM+wOleZbkhUrhKG6ctFR2W6mur8V1D/LZGnugVB
gASnV9xJzvgOEsfEt+BDInrVa3foKprI0vqEhg2qGw27kqUgbWO4pyK6tr6LsyCucyRdYm0A4oj/
SNS6CoY96za3yqcOmhVSU5sFTkz49q7FjdyjYC9Pus7M/AwtYx3kRju9XuAeSddTxAs1klU5GV1w
ehW9OHgBnGUAV271ijZ6GgH25F8RBnXPDQkEd96o+7YY+HrytZIfZDsp1Xlf8LMKROL3VRwk/qHd
iitcovj/Fh9H1VGa7By8cS5jNQsSKsBaBfuE5Iz6LWF2qRELXiuuU1+r8OORcZZy+0TZ1RduF6rP
koW25HaJydJSNggEjb9TuuAEIeiXOARDg/EYui2Q43xHcSkN1JelN4nze+0e9RjDS0FlREmqqBFz
26bES2BJ8ho6X6pU/nDvautk8xZPPh3R6T3tkOMTKv/Qb2BuNErs7Ff5qryxMOzwOV+Os6/DSErq
VA1pwZzC5jtARwpv72OXGmlhrjDCIw4jj1DGHW+i8J3SFWyYN8UmMWHtZfWq7VKtqnd6QxXJxGh4
1ID0xvIYDrgp72R7Ni8ykMwv5igb8pJ+5f5guYZ15XcA2SAdi6I1kxMXJGAGr6dYOXHf2TTfRQta
0Z/t/pbzDzxZhUX9DpO9MVq9tQR9vpv9UQ5BhmT66Xehj34DmPdSRZbP6xFfw/e9YqSmauXJF7L4
Vm0EIrKmGWFjgNONtYiRc16AHCjg8xSsOgxRsFnmSdiA4n/bprYZtX+OP5xo2KpffzyZIWku2CA9
RDeB/Sgnv8EAowwK8LOhZK+n0kTGby8a9iI9EJby87RCVV6+kP+QMbY6J88MY17em9VX/x2+fOy9
S94Bav+g67FEm+XqwakVAe9fRXWG6+2rLS1v9DJmI3oByw3yC9zJZvvZkakiUGBqRHH1ehxn0iwe
Ii2dYj5argb49PFX3cIeyu2I7JeR4PT+5uSxw9DBlx7pdBQhMZfXyIAElmEYpoaZzyi0xanMU68q
jv8vyIsWxKKLLD257wQA0hFDrs39Nl4ZjsdZ2e/5TnxwvWWif1AsJ3kuAhcKVZ4RbUceWZyqIH5d
j1c+WKLnJ4Vb+ORx6RtH4EHmU+2mj9BvnVqCBna069TvhICDGHMrR9sL81YRGmSi8Isnz0tE823o
HiNbuCXGLg8/TIpojSlvQyByHSN70pMoloHIP5Lfplh6gWxq5ZZqQ9O+9ImiEFy+8K/KNy50/o9I
tHTeahTrYJtn7YmV2BlqM48adCVhEB44WvXB6B1g557akamUiXsMA7d2X7SCZUfXYvRqeFnSZsro
iCywN55yU94OVhqj6HETov2utJdH5QV2FFvSDsh2gM7MC8laGjBbJMAheVlpIx7/QYuLTorfSyJf
rxXpkwUIJgIf1PzhgYzuepUsH6LBIPCQ2VjU/cRyk/+WswsbAizlDEDRh9bJnvmzYXHJNxB5B9Oj
tQ7Os4LnUVJTmEBzcrkBV94/6HIkYVaAb6WTj6n3sq7lbjF4wd3/yLvusVVYKMm+0sUP6Zd6rG/9
n/BB3Dn81lu8YMiKkkE5DOBo6nLL8V45PYVqOc5a1ZoWHXq3EZPJapOTDP/wZ0+CV8gUrptDRswf
eonYkLUWnZ2r7GVFsgIGIshtivud5AWE5EfOU2xUNZyzyj2/fOqdPpjUwnudKfVzH1DrMGuhK772
i/mlEX5bsCMdQF4Wll5vchjAo8Dmp1TWP3WuSqXpgsEP+I0OgtiIowY6Yi6+gHHtxJo4BW5pPE3F
ZeSUkkrcp+fhgxPgrCGdz62fe5hUgfZQMDchJaVNs+XIZjOHhz8kDM+KawhDPoAuHfzNU+faaVHo
tfmVE6zailldqs36cJdprMKooSN1EiTBZN8YK7506m0qMuehN8ABMt7ac18NTd3j/8bmoQPB8/Gr
FjaOWA4xCTFQnV3hTn+2euCDW+pTb4cQgzpLlQWSW5Xh5hQHdN8iZ6Bj785rXuehbdWhpLU223Qx
WRKkAZWiodb8dsQfSsT1ONqs7sbmaxC2zKaFfWiIrh92GSShfELyLKWAXE/8kC1wPdXz4H5rsKMB
ZZGoBoUacTLnisxhSzceiyLxn+k0vJwDZLUFDEtLdhaxIe9lZrDzoc5AJ2m9Wyeib9XI7+r9I/oc
JO/7Oxc97AQCOWVx1rVlv3wZYYArboA2Pqz82XluCnkJYNDV6WbJsxgG+wQCPmwYW2PEY9udtt3E
dJy5AcNc7G5W+UsHSyV4KfoZCwkSK6wxCGN5a/BVhhP46ffwbLfNDZEA03j32H2ArPVrIR1VEuyl
Gk0EdjsbUUuKmVG00gau+UvF7a1/Ga7F1IV5xptOM15Of/7Ro28/EqFQ5QPwXM1Qljw94xhprhXA
dxgU7IGTPtB/H4d6GZv2C9lpP2ZZ9aakCdiU+vgz1dUpXwVQiM0oocb8wdFb2tNvDXz/ITfT/Hcy
E/hEbKfG8xC1iliOLW6fPsCqvMcdWqdw6M6iTAROoCwCeLU7Z8bf1XNkjku0B9fuywTLapmnF6xu
kt4oLLsrRNHJW6iP+7f8Gl1CbgbxqVx4aRTg7iTpTGepcup3rJDKBP9Vul3g2RAce0ttu/Vey1dq
uhYBzqf2/tEHuvzBVY2xkKs+BNOY2ljprwQyPTRc7k7ndZJz8SXqOoCp0cEs4rO45GQ+Vc0tWcQN
eX6zV9q6innILimaPDRHghqADdojYppg9aM/Srbn2vQWLDjIdKXxmWSoYntxn1nu14uZap3nR3GZ
vajYQE3YC7MLJ7SRGENogo2IQ2aVdeE83fZzVAHmabMi92AZNULUlGCWwLV1x7l9Puc2lFHVwq3X
LsG9vCxlmYYUETYL7ygC0u7jIFXchp0RJbwgtwH01hhEHQ4ekdDKGExuAlSoLoSBdGC8f9+SGBDp
q+McGkBJqhf8wk2fmnyvZeN8slRADTZhD2hFY2nHO8oZRw4Pl9yeuewcav+Q3ohvjVOG657vEsnZ
yarYBI6HXMJ9V4rXKZTJGZE5nOihZKOnQ0w7+A4AxLruTu0eFQGv/DHa+3LWGCx2th3qmKU9Cffi
gSNsHxCTeOUO+XNGr7JKXbO5QoRurGkrC6zd4xzByFRLIXaYJ559AGi7n8UwOiIYtE32bJwSeT6c
lzwxWo+Gebo2JYmLLfCTg6ZRGbppO52oNk1P6GvT8RVlzLYXLN3tlGpbhst8neeGxVv8DB2dzRSD
oYePMJU1kWSxiPz9rJ4TG0vej1x05BVUAIjUIaVcOUuuWW6LJeQ7osusH6XpgXyi0Mn/9wFwhdnx
I01BBFfpHIbaianYMDJzEZbf4FXUvNlP4JnVqzoRYIx2rlgsM4cCPgGkLvxK4ZG5NAmPCsj+k9yM
8qHLmL7cc9Vfq/ISg3cVhZ76em38UEyWK+S35B4zCPRjBOgOfbNoAFSfJ5Qs3tU6cwpTboBnew6q
zWtpJSMkeBD9dJLtU3lbCo8uUfDnHSUo6o9CdSn03SXgOGChpytpSWkTWo/dmhLpll3IaQDiaCVU
dZPrt1ui9gZB1pc4XMEqwnQ2G1gBQxFsfW6SdTaNjPlsoBK/l/jxELumOH8Msu5yWvqjd2a6skFp
Z2T5clCBC5t24ADNf6CK4b1Tm8BqUvfIDcQxzSgPXojH1P39k+4CJt2ivTwnXxCcW2i4RD9fLPkb
ZRcmRVyxoBOXFP1v4UGwabGsKPhSa29IGTuu+2VBVycKuwV3aVDlq9OV8CWXjg2EoBuMMW2N963f
vQy+Uag34loYourh4V4qEyr6GgMLXFYm5xu6p5Ob0wZt/zWLHDWjUbPcEVveMN0Cd0eDP2du7izL
t+KbXV/+yzvHoSojjUJTV+qsNfJQuc+0gqtZ9gHRUtYqLowhMN0zWDg5ugtQNuw6PLXsgswozioG
G6dG59xSV685v0hlo7SUG68DnAYX+XYR4TREFbLBuUlK+qCpNvEsaYwd7J5D+sfbLjnf4ekgh10v
DRTV123I5ZRL89whJrWhapZ+K9uGmorwYZAsVOhGN/wvZY+Q0wsOGPkf7TSQt/8Uk+qP3CaSOkO/
NVVJQWZQDuo+2UDPQ1CNHuEOgznFadK5LTTDG9ugxUrSYc5O/gi1wVf+w89S3vp4orS8TQkpOp3A
bax4sHbf1n2PyCvifAjh0G77jQ1x9nVwa205X7RhvOxZFsw2qJc189O4EHOuADpAuWy9QShGqzyG
oPeFVj+9YJjsecgxHdoBp8aUTTjV8T3nyZGxmvEXoP8RB7gOtjjg5855JVcyj7r+Dh5CJV9sP4NW
icu7c8t97EPOwHblPHz+jzSPtR5d9CYujm9V7SOP8StgpRvy4kKqhO1cPzbwAVZRPCdQq+MQnxiZ
4caBkd3ozYtG4MGJzY8AvpBa7GnCu2RTY99gLNx/tyC0CiMYAYSXAB4zA83mSLWVd5PsEHIvhgz+
9h0GrkomhqcVjZpJLoDH3AAYKXesLdUbKD6+HLt118Ql9FRdL0K03JAb2CzHfzlD4NZitxjWCQ8l
GU1ED0bUmDtuC5rXFcdFM9aEonGkvDV5qQ6EazWXWR+aFVninVfAgCTyX2hAHewte6413etbCT20
A0P5pDB7QHQT3M5k9fRRjnoe46wSbZKR61HcZQ40G+rPPFEI1WW67TGZE0TylBFBtt6mdqWOxkI4
E005UiaxbNiSdF/LYDBuxCgmD0pGu4ojjuxv9yAA53bB8zmJpcir5gZKN5noAg3lPQLLkt5fKaTM
x4k6C6QnqoPvrN0SJcyjkbQAiXdD69YO4Udpx1WMxEKgkePAByFm9s2XswetEHD/vQbOzq7i3tFr
65eLUZx8z1XMLF1F9L1peXjOUADIgXmOkiydqklVF7ZGXnn8doB/dlE9somuAtuOqn9J6AWkWaTw
IISw0CrlKNkJZso6Y3e+SmF1S9+bWmuMKZb1tnWZMqrq2SShaZH6R9mrQ2F6DO6d3f0+nTCbMVdz
mvCbbPhroflpuxqDHb1/e6BVTRbTOSd8kCGmyFv64gLdW3jznsTsQuVIVEg9DW9+MryvtMC8ng70
l2hRmwrNeY51vv3/3aGDeH1T19fwAeGO9XwnxAwxb5O6ZrLpQZMBqz+x0vfXufdxcV+UvDpA3qrM
GJG7fJYkTterm+7S9FxG0WisfziBPxokF2gLsNBWEPaxWCwHhgv8UGYhvvq4sMA/anjU+IRHi2qz
1Smz3diwbRLNjty5xF6Wh0joxGF5GFkniaK7MXBFHS+kzm7Ea2hFmIaYWwo/mM1n9ap4TgI7n0FO
2gpiyHUokapZqNEW0o6bbAGUJClsKlb1GKeOEziDxkRTdgjcZ1iEfjSFToJ6E5OFgDkz/FrVocCL
lylla0tQeRxEfbW0046VrhM75A92lDUFxnMSBR3LElzuBUnuA5E5VuEssXmjhXa/Jko0mYxVjYzH
KLIymqdd2rUgpDubjzqvws4lAI2PiGNvydJ9TcC+vS6gmMuXCdqtXbd3qiyechk9JiVQjGhdoKJN
UtDpKjZVwJxcNcrvX9NSa87tDzJmriDntYXPGd0NyeDKK9Ibou1+vFi3MYu8W/ki+UUdURsX6W+J
yxU2QhrKT7sRHVCcJGzaDl88WYZOHQsq5rf5i+xqtA8N+1O4MugXZjwlKzXRJiZIBq1CHZ5tw7GU
YWmqAKeEMabrE7SCcbU3dVSwUSkHnJrdp2G6kXdSjZXj9mXN/dE+iUbioYK1fFm/sI2UvdI3vGW/
V7rhN0HV5wn8VdBvn9m4xax5vrNL02gPa8FI1jlt8ShW4mBC8Mj607U1r4nWxWSMlEEbkvLiPUC5
WEXfdluSG4H4/W5eJx+9WUI=
`pragma protect end_protected
