`ifndef DMA_DEFINES_VH
`define DMA_DEFINES_VH


`endif

